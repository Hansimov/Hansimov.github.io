MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       �+K�J{�J{�J{o��J{ߌ�J{ߌ�J{;E&�J{�Jz�J{ߌ�J{ߌ�J{ߌ�J{Rich�J{                        PE  L K?eL        � !  �  �      ��     �                         `                              p� J   � (                            0 �!                                  p� @            �                            .text   5�     �                   `.rdata  �3   �  @   �             @  @.data   �4   �      �             @  �.reloc  �-   0  0                @  B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        U��`V��H�QV�ҡ`�H�U�AVR�Ѓ���^]� U��`V��H�QV�ҡ`�U�H�E�IRj�PV�у���^]� ����������U��`�H�U�I(��VWR�E�P�ы`�u���B�HV�ы`�B�HVW�ы`�B�P�M�Q�҃�_��^��]���U��`�H�A�U���R�Ћ`�Q�Jj j��E�hp�P�эU�R��  �`�H�A�U�R�Ѓ���]��������������U��`�H�A�U���R�Ћ`�Q�Jj j��E�h��P�эU�R�  �`�H�A�U�R�Ћ`�Q�J�E�P�ы`�B�Pj j��M�h��Q�ҍE�P�N  �`�Q�J�E�P�ы`�B�P�M�Q�ҡ`�H�Aj j��U�hp�R�ЍM���LQ�  �`�B�P�M�Q�҃���]������������U��MW�};�u3�_]ËE�U��PS�X;�u[3�_]�V�0;�t;�u�p;�tk;�tg�p;�t;�u;�tV;�tR;�t;�u;�t-;�t);�t;�uI�;�t;�u?�M�1�P�E^[��   _]Ë�U�
�@�M^[��   _]Ë�M��P�E�^[�   _]��������������U���T�`�HH���   SVW�}h�  W�ҋ�`�HH���   h�  W�u��҃��ωE���/  ���؉]���  ���BT  ����  �`�HH��p  j h�  W�҉E�`�HH��p  j h�  W�҃��E�P�M�Q���3�W�ˉu�u���T  ��t>�d$ �EԋM؃�;��I ���u����E��;�~�U�R�E�PW���T  ��uɉu�M�]������U��P�U��P�@�U��U����E��
��P�M��H�U��P�MĉU�3�3�3��D��;E�u��u	�   ����   �E�;E�u��u	�   ����   �E�;E�u��u	�   ����   �E�;E�u��u	�   ����   �E�����|��ɉ]��q  ���i  �} �S  �M��S7  �u�E�M�j VPQ�M��m7  �U��   ;��]��U�|p�E�M�PQS�M���7  �����tU�M�V�u��R  �Ǚ�}��t	�M�V�$S  �M��U�R�U�E�PQSVR���������t�]�;]�u�E�;E�t��;}�~��u���}��]܉}��]��E�    |r�d$ �M�QSW�M��B7  �����tY�M�V�u��/R  �E��}��t	�M�V�R  �M�U�R�E�PSWVQ�W�������t�}�;}��]�u;]�t�E��;E�E�~��`���   �M�Pj j��j �#  ���M��6  _^�   [��]�_^3�[��]��������������������U��E�� t"��t-�  t3�]ùh��  �����]ø   ]�������������U���$Vh'  ��  ��`�H�A�U�R�Ћ`�Q�J�E�PV��h`�jjh�j�]  ���� ��t���T  ���3��`�B�P�M�Q�ҡ`�H�Aj j��U�hP�R�Ѓ��M�Q�M��A�  � V�U�RPj ��Phٞ �
V  ���M����=�  �`�Q�J�E�P�ы`�B�P�M�Q�҃���^��]����������������U��`�H�Q��@V�uV�ҡ`�H�Qj j�h(�V�ҍE�jP�����`�QVP�B�Ћ`�Q�J�E�P�ы`�B�P�M�Q�ҡ`�H�Aj j��U�h��R�ЍM�j Q�]�����DP�U�R�E�VP�[
  ��P�M�Q�N
  �`�J�QVP�ҡ`�H�A�U�R�Ћ`�Q�J�E�P�ы`�B�P�M�Q�ҡ`�H�A�U�R�Ћ`�Q�J�E�P�ы`�B�Pj j��M�h��Q�ҍE�j P������@P�M�Q�U�VR�	  ��P�E�P�	  �`�QVP�B�Ћ`�Q�J�E�P�ы`�B�P�M�Q�ҡ`�H�A�U�R�Ћ`�Q�J�E�P�у�$��^��]�U��`�H�A�U���`R�Ћ`�Q�Jj j��E�h(�P�эU�R�����`�Q�R�M�QP�ҡ`�H�A�U�R�Ћ`�Q�J�E�P�ы`�B�Pj j��M�h�Q�ҡ`�H�A�U�R�Ћ`�Q�Jj j��E�h�P�ы`�B�P�MЃ�LQ�ҡ`�H�I�U�R�E�P�ы`�B���MЋP<�ҋ`�Q�RLj�j��MQP�M��ҡ`�H�A�U�R�Ћ`�Q�R�E�P�M�Q�ҡ`�P�B<���M��Ћ`�Q�RLj�j��M�QP�M��ҡ`�H�A�U�R�Ћ`�Q�R�E�P�M�Q�ҡ`�P�B<���M��Ћ`�Q�RLj�j��M�QP�M��ҍE�P��  �`�Q�J�E�P�ы`�B�P�M�Q�ҡ`�H�A�U�R�Ћ`�Q�J�E�P�ы`�B�P�M�Q�҃��} tH�`�H�A�U�R�Ћ`�Q�Jj j��E�h�P�эU�R�h  �`�H�A�U�R���H�`�Q�J�E�P�ы`�B�Pj j��M�h��Q�ҍE�P�  �`�Q�J�E�P�ы`�B�P�M���Q�ҡ`�H�A�UR�Ѓ���]�U���$Vh'  ���  ��`�H�A�U�R�Ћ`�Q�J�E�PV��h`�jfh�j�vW  ���� ��t���vN  �0��3��`�B�P�M�Q�ҡ`�H�Aj j��U�h�R�Ѓ��M�Q�M���  � V�U�RPj ��Ph؞ �jP  ���M�����  �`�Q�J�E�P�ы`�B�P�M�Q�҃���^��]����������������VW���������Ph'  ��  ���`�H�Q����V�ҡ`�H�QVW�҃������������Ph'  調  ���`�H�Q����V�ҡ`�H�QVW�҃�����������_�   ^���������������U���Vhٞ ���  ����tF�`h���h  �j jj
j�E��  �E�    �Qj�ȋ��   h�  ��P�M�Q���pa  �   ^��]�������U��� SVW��� �  h'  ���Ծ  �ء`�H�A�U�R�Ћ`�Q�J�E�PS�у��U�R���_  �`�H�A�U�R�Ћ`�Q�Jj j��E�h(�P�у�j �U�Rj jj?j ���,}  �`�H�A�U�R�Ѓ�jjjj����}  jj���^}  �`�Q�J�E�P�ы`�Bj j�h(��M��PQ�҃�j �E�Pj jj j ���|  �`�Q�J�E�P�у�j j j j ���}  jj����|  j �U�Rj j jh�  ���t  j jFjh�  ��� w  ���|  jj ���~r  j����}  ���~|  h���h  �j jj
jj�E�P���E��  �E�    �_  �`�Q�J�E�P�у���_^[��]����U���V�qV�E�P�E��  �E�    ��e  �M��6�  �`��Q�R4Ph�  �M���j�E�Phٞ �]
  ���M��b�  3�^��]������������U���VW�}���~�  ������   �`���   �Bh�  ���Ѕ���   �M���  hk/  �E���E�    �  ����urh�?  �t  ����uah�/  �c  ����tPjjV���������t?j j j j�j��M��)�  �}� t'����  Vj+���B�  �M�j QV����������  �M��ă  _�   ^��]� ������̸   @� ��������U��V��蕃  �Et	V�Q  ����^]� ���������������U��VW�}���Q�  ������   �`���   �Bh�  ���Ѕ�tihk/  �r  ����uXh�?  �a  ����uGh�/  �P  ����t6jjV���������t%����  Vj+���G�  j jV����������  _�   ^]� ��������U��V���H  �Et	V�P  ����^]� ���������������U��`�H�QV�uV�ҡ`�H�U�AVR�Ћ`�Q�B<�����Ћ`�Q�M�RLj�j�QP���ҋ�^]���������U��E�`� ]��U��`�P8�EPQ�JD�у�]� ���̡`�H8�Q<�����U��`�H8�A@V�u�R�Ѓ��    ^]�������������̡`�H8�������U��`�H8�AV�u�R�Ѓ��    ^]��������������U��`�P8�EP�EP�EPQ�J�у�]� ������������U��`�P8�EP�EPQ�J�у�]� �`�P8�BQ�Ѓ����������������U��`�P8�EPQ�J �у�]� ����U��`�P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U��`�P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U��`�P8�EP�EPQ�J(�у�]� U��`�P8�EP�EP�EPQ�J,�у�]� ������������U��`�P8�EP�EP�EPQ�J�у�]� ������������U��`�P8�EP�EP�EP�EP�EPQ�J�у�]� ����U��`�P8�EP�EPQ�J0�у�]� U��`�P8�EP�EP�EPQ�J4�у�]� ������������U��`�P8�EPQ�J8�у�]� ����U��`�H��x  ]��������������U��`�H��|  ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H�A,]�����������������U��`�H�QV�uV�ҡ`�H�Q8V�҃���^]�����̡`�H�Q<�����U��`�H�I@]����������������̡`�H�QD����̡`�H�QH�����U��`�H�AL]�����������������U��`�H�IP]�����������������U��`�H��<  ]��������������U��`�H��,  ]��������������U��`�H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡`�H���   ��`�H���  ��U��`�H�U�ER�UP�ER�UP���   Rh�.  �Ѓ�]����������������U��`�H�A]�����������������U��`�H��\  ]��������������U��`�H�AT]�����������������U��`�H�AX]�����������������U��`�H�A\]����������������̡`�H�Q`����̡`�H�Qd����̡`�H�Qh�����U��`�H�Al]�����������������U��`�H�Ap]�����������������U��`�H�At]�����������������U��`�H��D  ]��������������U��`�H��  ]��������������U��`�H�Ix]�����������������U��`�H��@  ]��������������U��V�u����  �`�H�U�A|VR�Ѓ���^]���������U��`�H���   ]��������������U��`�H��h  ]��������������U��`�H��d  ]��������������U��`�H���  ]�������������̡`�H���   ��U��`�H��l  ]��������������U��`�H��   ]��������������U��`�H��  ]��������������U��V�u����  �`�H���   V�҃���^]���������̡`�H��`  ��U��`�H��  ]��������������U��`�H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U��`�H���  ]��������������U��U�E�`�H�E���   R���\$�E�$P�у�]�U��`�H���   ]��������������U��`�H���   ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H���   ]��������������U��`�H���   ]��������������U��`�H���   ]��������������U��`�H���   ]��������������U��`�H���   ]��������������U��`�H���   ]��������������U��`�P���E�P�E�P�E�PQ���   �у����#E���]����������������U��`�P���E�P�E�P�E�PQ���   �у����#E���]����������������U��`�P���E�P�E�P�E�PQ���   �у����#E���]����������������U��`�H��8  ]��������������U��V�u(V�u$�E�@�`�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@�`�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��`�P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U��`�P0�EP�EP�EP�EPQ���   �у�]� ����̡`�P0���   Q�Ѓ�������������U��`�P0�EP�EPQ���   �у�]� �������������U��`�P0�EP�EP�EP�EPQ���   �у�]� ����̡`�P0���   Q�Ѓ������������̡`�H0���   ��U��`�H0���   V�u�R�Ѓ��    ^]�����������U��`�H��H  ]��������������U��`�H��T  ]�������������̡`�H��p  ��`�H���  ��U��`�H���  ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H�U�E��X  ��VR�UPR�E�P�ыu�    �F    �`���   �Qj PV�ҡ`���   ��U�R�Ѓ� ��^��]��������U���$Vj hLGOg�M����  P�E�hicMCP�k������M�� �  �`���   �JT�E�P�у���u(�u��蚺  �`���   ��M�Q�҃���^��]á`���   �AT�U�R�Ћu��P��蚺  �`���   �
�E�P�у���^��]�������������U��`�H��  ]��������������U��`�H��\  ]��������������U��`�H�U��t  ��V�uVR�E�P�у����s�  �M���  ��^��]�����U��`�H�U���  ��VWR�E�P�ы`�u���B�HV�ы`�B�HVW�ы`�B�P�M�Q�҃�_��^��]����������������U��`�H�U���  ��VWR�E�P�ы`�u���B�HV�ы`�B�HVW�ы`�B�P�M�Q�҃�_��^��]����������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H�U�E��VWj R�UP�ERP��t  �U�R�Ћ`�Q�u���BV�Ћ`�Q�BVW�Ћ`�Q�J�E�P�у�(_��^��]��U��`�H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    �`���   j P�BV�Ћ`���   �
�E�P�у�$��^��]���U��`�H��8  ]��������������U���  ���3ŉE��M�EPQ������h   R�Ͽ ����|	=�  |#��`�H��0  h0�hF  �҃��E� �`�H��4  ������Rht��ЋM�3̓��w� ��]�������U��`�H��  ��V�U�WR�Ћ`�Q�u���BV�Ћ`�Q�BVW�Ћ`�Q�J�E�P�у�_��^��]����U��`�H��  ��V�U�WR�Ћ`�Q�u���BV�Ћ`�Q�BVW�Ћ`�Q�J�E�P�у�_��^��]����U��`�H��p  ��$�҅�trh���M��ٵ  �`�P�E�R4Ph���M��ҡ`�P�E�R4Ph���M���j �E�P�M�hicMCQ�����`���   ��M�Q�҃��M�贵  ��]�U��`�H��p  ��$V�҅�u�`�H�u�QV�҃���^��]�Wh!���M��,�  �`�P�E�R4Ph!���M���j �E�P�M�hicMCQ�����`���   �QHP�ҋu���`�H�QV�ҡ`�H�QVW�ҡ`���   ��U�R�Ѓ�$�M���  _��^��]������U��`�H��p  ��$V�҅�u�`�H�u�QV�҃���^��]�Wh����M��\�  �`�P�E�R4Ph����M���j �E�P�M�hicMCQ�����`���   �QHP�ҋu���`�H�QV�ҡ`�H�QVW�ҡ`���   ��U�R�Ѓ�$�M���  _��^��]������U��`�H��p  ��$�҅�u��]�Vh#���M�褳  �`�P�E�R4Ph#���M���j �E�P�M�hicMCQ������`���   �Q8P�ҋ�`���   ��U�R�Ѓ��M�腳  ��^��]���������������U��`�H��p  ��$�҅�u��]�Vhs���M���  �`�P�E�R4Phs���M���j �E�P�M�hicMCQ�W����`���   �Q8P�ҋ�`���   ��U�R�Ѓ��M���  ��^��]���������������U��`�H���  ]��������������U��`�H��@  ]��������������U��`�H���  ]��������������U��V�u���t�`�QP��D  �Ѓ��    ^]������U��`�H��H  ]��������������U��`�H��L  ]��������������U��`�H��P  ]��������������U��`�H��T  ]��������������U��`�H��X  ]��������������U��`�H��\  ]�������������̡`�H��d  ��U��`�H��h  ]��������������U��`�H��l  ]�������������̡`�H���  ��U��`�H�U���  ��VR�E�P�ыu��P���Ӱ  �M���  ��^��]�����U��`�H���  ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H���  ]��������������U��`�H��$  ]��������������U��`�H��(  ]��������������U��`�H��,  ]�������������̡`�H��0  ��`�H��<  ��U��`�H���  ]�������������̡`�H���  ��U��`�H���  ]������������������������������U��`�H��  ]�������������̡`�H��P  ��`���   ���   ��Q��Y��������U��`�H�A�U��� R�Ћ`�Q�Jj j��E�hx�P�ыUR�E�P�M�Q�-����`�B�P�M�Q�ҡ`�H�A�U�R�Ћ`�Q�J�E�P�у�,��]��U��`�E�PH�B���$Q�Ѓ�]� ���������������U��`�PH�EPQ���   �у�]� �U��`�PH�EPQ���  �у�]� �U��`�PH�EPQ���  �у�]� �U��`�PH�EP�EPQ��  �у�]� �������������U��`�PH�EP�EPQ��  �у�]� ������������̡`�PH���  Q�Ѓ�������������U��`�PH�EPQ���  �у�]� ̡`�PH���   j Q�Ѓ�����������U��`�PH�EPj Q���   �у�]� ��������������̡`�PH���   jQ�Ѓ�����������U��`�PH�EPjQ���   �у�]� ��������������̡`�PH���   jQ�Ѓ����������U��`�PH�EPjQ���   �у�]� ���������������U��`�PH�EP�EPQ���   �у�]� �������������U��`�PH�EP�EPQ���   �у�]� ������������̡`�PH���   Q�Ѓ�������������U��`�PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP�����  ������t�E�`�QH���   PVW�у���_^]� �����U��EVW���MPQ���  ������t�M�`�BH���   QVW�҃���_^]� ̡`�PH���   Q�Ѓ������������̡`�PH���   Q�Ѓ�������������U��`�PH�EPQ���   �у�]� �U��`�PH�EPQ���   �у�]� �U��`�PH�EP�EPQ��8  �у�]� �������������U��`�PH�EP�EPQ��   �у�]� ������������̡`�PH���  Q�Ѓ������������̡`�PH���  Q�Ѓ������������̡`�PH���  Q�Ѓ������������̡`�PH��  Q�Ѓ������������̡`�PH��  Q�Ѓ�������������U��`�PH�EP�EPQ��  �у�]� �������������U��`�PH�EP�EP�EPQ��   �у�]� ���������U��`�PH�EP�EP�EP�EPQ��|  �у�]� �����U��`�PH�EPQ��  �у�]� ̡`�PH��T  Q�Ѓ�������������U��`�PH�EP�EPQ��  �у�]� �������������U��`�PH�EPQ��8  �у�]� �U��`�PH�EPQ��<  �у�]� �U��`�PH�EPQ��@  �у�]� �U��`�PH�EP�EP�EPQ��D  �у�]� ��������̡`�PH��L  Q��Y��������������U��`�PH�EPQ��H  �у�]� ̡`V��H@�Q,WV�ҋ`�Q��j �ȋ��   h�  �Ћ`�QH�����   h�  V�Ѓ���
��t_3�^Ë�_^�̡`�P@�B,Q�Ћ`�Q��j �ȋ��   h�  �������U��`�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U��`�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U��`�PH�EP�EP�EPQ��   �у�]� ��������̡`�HH��  ��U��`�HH��  ]��������������U��`�E�PH��$  ���$Q�Ѓ�]� �����������̡`�PH��(  Q�Ѓ�������������U��`�PH�EP�EPQ��,  �у�]� �������������U��`�E�PH�EP�E���$PQ��0  �у�]� ���̡`�PH���  Q�Ѓ������������̡`�PH��4  Q�Ѓ������������̋��     �������̡`�PH���|  jP�у���������U��`�UV��HH��x  R��3Ƀ������^��]� ��̡`�PH���|  j P�у��������̡`�PH��P  Q�Ѓ������������̡`�PH��T  Q�Ѓ������������̡`�PH��X  Q�Ѓ�������������U��`�PH��Q��\  �E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����̡`�PH��`  Q�Ѓ�������������U��`�PH�EPQ��d  �у�]� �U��`�E�PH��h  ���$Q�Ѓ�]� ������������U��`�E�PH��t  ���$Q�Ѓ�]� ������������U��`�E�PH��l  ���$Q�Ѓ�]� ������������U��`�PH�EPQ��p  �у�]� �U��`�PH�EP�EP�EP�EPQ���  �у�]� �����U��`�PH�EP�EP�EP�EP�EP�EPQ���  �у�]� �������������U��`�E�HH�U �ER�UP�E���$R�UP���   R�Ѓ�]������������U��U�E�`�HH�E���   R�U���$P�ERP�у�]����������������U���E�M����L� �M;�|�M;�~��]�����������U��`�PH�E���   Q�MPQ�҃�]� ������������̡`�PH���   Q��Y�������������̡`�PH���   Q�Ѓ������������̡`�PH���   Q��Y��������������U��`�PH�EP�EPQ���   �у�]� �������������U��`�PH�EP�EP�EP�EP�EPQ���  �у�]� ̡`�PH��t  Q��Y�������������̋�� ���@    �����`�Pl�A�JP��Y��������U��`V��Hl�V�AR�ЋE����u
�   ^]� �`�Ql�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uË`�QlP�B�Ѓ�������U��`�Pl�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U��U�E�`�HH�ER�U���$P���  R�Ѓ�]����U��`�HH���  ]��������������U��`�HH���  ]��������������U��U0�E(�`�HH�E$R�U ���$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�,]������������U��`�HH���  ]��������������U��`�E�PH�EP���$Q���  �у�]� ��������U���SV���  �؅ۉ]���   �} ��   �`�HH��p  j h�  V�҃����E�u
^��[��]� �MW3��}��   ����   �]��I �E�P�M�Q�MW��  ��tc�u�;u�[�I ������u�E�������L�;Ht-�`�Bl�S�@����QR�ЋD������t	�M�P��  ��;u�~��}��M���}��  ;��r����]�_^��[��]� ^3�[��]� ����������U����`SV�ًHH��p  j h�  S�]��ҋ�����u
^3�[��]� �E��u�`�HH���  �'��u�`�HH���  ���uš`�HH���  S�ҋȃ��ɉEt�W�T  �`�HH���   h�  S3��҃����  ���_�u����    �`�Hl�U�B�IWP�ы�������   �`�F�J\�UP�A,R�Ѓ���t�K�Q�M�u  �`�F�J\�UP�A,R�Ѓ���t�K�Q�M�L  �E��;Pt&�F�`�Q\�J,P�EP�у���t	�MS�  �`�v�B\�M�P,VQ�҃���t�M�CP��  �`�QH�E����   �E�h�  P�����у�;�����_^�   [��]� ������U��`�HH���   ]�������������̡`�PH���   Q��Y��������������U��`�HH���  ]��������������U��`��P���   V�uW�}���$V�����E������At���E������z����؋`�Q�B,���$V����_^]����������������U���0��`�U�V�u�U��]�W�P�}���   �E�PV�M�Q����� �@�@�E�����E��Au�����������z���������������z�����������Au������������z)���١`�]��ɋ��]��]��P�RH�E�PV��_^��]���������Au������������������U��`�HH�]��U��`�H@�AV�u�R�Ѓ��    ^]�������������̡`�HH�h�  �҃�������������U��`�H@�AV�u�R�Ѓ��    ^]��������������U��`�HH�Vh  �ҋ�������   �EPh�  � �  ����t]�`�QHj P���   V�ЋMQh(  ���  ����t3�`�JH���   j PV�ҡ`���   �B��j j���Ћ�^]á`�H@�QV�҃�3�^]�������U��`�H@�AV�u�R�Ѓ��    ^]��������������U��`�HH�Vh�  �ҋ�����u^]á`�HH�U�E��  RPV�у���u�`�B@�HV�у�3���^]�������U��`�H@�AV�u�R�Ѓ��    ^]��������������U��`�HH�I]�����������������U��`�H@�AV�u�R�Ѓ��    ^]��������������U��`�PH�EPQ���  �у�]� �U��`�PH�EPQ���  �у�]� ̡`�PH���  Q�Ѓ�������������U��`�HH���  ]��������������U��`�E�HH�U0�E,R�U(P�E$R�U P�ER�U���\$�E�$P��P  R�Ѓ�,]������������̡`�PH���  Q�Ѓ�������������U��`�PH�EP�EPQ���  �у�]� ������������̡`�PH��  Q�Ѓ�������������U��`�PH�EP�EP�EPQ���  �у�]� ��������̡`�PH���  Q�Ѓ������������̡`�PH���  Q�Ѓ�������������U��`�PH�EPQ��  �у�]� �U��`�PH�EPQ��  �у�]� ̋������������������������������̡`�HH���  ��U��`�HH���  ]��������������U��`�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ���������U��`�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ��������̡`�PH��,  Q�Ѓ�������������U��`�PH�EPQ��X  �у�]� ̡`�PH��\  Q�Ѓ�������������U��`�HH��0  ]��������������U��`��W���HH���   j h�  W�҃��} u�   _��]� Vh�  ��  ��������   �`�HH���   j VW�҃��M�胓  �`�P�E�R0Ph�  �M����E�`�P�B,���$h�  �M��Ћ`�Q@�J(j �E�PV�у��M�茓  ^�   _��]� ^3�_��]� �����U��S�]�; VW��u7�`�U�HH���   RW�Ѓ���u�`�QH���   jW�Ѓ���t�   �����   �`�QH���   W�Ѓ��} u(�`�E�QH�M���  P�ESQ�MPQW�҃��B�u��t;�`�U�HH�ER�USP���  VRW�Ћ`���   �B(�����Ћ���uŃ; u�`�QH���   W�Ѓ���t3���   ���Wu1�`�QH���   �Ћ`�E�QH���   PW�у�_^[]� �`�BH���   �у��} u0�`�M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� �`�QH�h  �Ћ؃���u_^[]� �`���   �u�Bx���Ћ`���   P�B|���Ѕ�tU�`�E�QH�MP�Ej Q���  VPW�у���t�`���   �ȋBHS�Ћ`���   �B(���Ћ���u�_^��[]� ��������������U��E��V��u�`�HH���  �'��u�`�HH���  ���u�`�HH���  V�҃���u3�^]� P�EP���>���^]� ���������U���D�`�HH���   S�]VWh�  S�ҋ�`�HH���   3�Wh�  S�u܉}��҃�;��E�}�}��}��p
  �`���   �B����=�  �`�  �QH���   Wh:  S�Ћ`�QH�E����   h�  S�Ћ`�QHW�����   h�  S�uԉ}��Ћ`�QH�E苂  S�Ћ`�QH�EЋ��  S�Ѓ�(���E��E����}   �M���M�MЅ�tMj�W���  ���t@�@�Ẽ|� �4�~����%�������;�u/�����  ;E�~�E؋���  E���E�;Pu�E���E��E���;}�|��}� tv�u�j S���x�  ����  �����  ��tV����  �}�;�uK�`�H���  �4�h����h�  V�҃����E��k  �M�PVP�z�  P�d ����}ܡ`�H���  �4�h����h�  V�҃����E��   �M�3�;�t;�tVQP��u ���E�;�~-�`�Qh����h�  P���   �Ѓ�;ǉE���  �`�E��QH��  j�PS�у�����  �u�;�tjS���Z�  ����  �����  �E���}�`�BH���   Wh�  S�у�3�9}ԉE�}���  �}���}ȋMЅ��p  �U�j�R���  ����\  �M̍@�|� ���]�~����%�������9E��  ����  �E�3�3�9C�E܉M���   ��I �����������t{�]��}������������ϋ9�<��}����҉��y�]��|��]������z�<��y�]��|��]������z�<��I�}��]������M��}ȃ��������M؃�;K�M��b������E��O  �+U�j��PR�M��c�  �M�v���E�3�+��U��E����	��$    ���E�;E���   �}� �U����E�t6�U�@�U�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�M��E�;]؍@�E��Ћ��P�Q�P�Q�P�Q�P�Q�@�A}c�UȋE�9�uX�ȋL�����������w4�$��f �U����4�"�M����t��U����t�
�M����t�M���;]�|��E�����;]؉M������U�;U��  �U�R�  �E�P�x  �M�Q�o  ��_^3�[��]Ë�M�3�;G�Å���   �E�v�ЋW��R�ы��Q�P�Q�P�Q�P�Q�P�I�H�O��I�M�ы�P�Q�P�Q���ۉP�Q�P�Q�P�I�H��@�E�ЋU�Lv�ʋ��P�Q�P�Q�P�Q�P�Q�@�At8�G�U�@�ʋU�Lv	�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��w��U��@�ʋU���v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��w��U����@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�7����t?�G�U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�w�����O�E�����;EԉE��}�������U�R�W  �E�P�N  ���$  ���   �B����=  �  �`�QH���   j h(  S�Ћ`�QH�����   h(  S�ЋЃ�3��҉U�~#���ǅ�t�|� t�4N��tN���;�|�u��u܋`�Q���  �4v�h����hK  V�Ѓ����E���   �M��t��tVQP��o ���u؋`�Q���  �h����hP  V�Ѓ����E�tP��t��tVWP�o ���M����+`�RH��PQ�E���   S�Ѓ���u�M�Q�  �U�R�  ��_^3�[��]á`�HH���   j h�  S�҉E��`�HH���   j h(  S��3�3���3�9]؉E��}ĉ]��N  �U���    �څ��+  ���E�    ��   �U�<��v��   ����U��:��\:�Y�\:�Y�\:׉Y�Z�Y�R�Q�U��\�E��Y�\�T���Y�Z�Y�Z�Y�Z�Y�R�]��Q�U�����������;�|��}ă|� �w   �U��Eԍ8�I�ʋU�v���A�B�A�B�A�B�A�B�I�J�E���ЋE���v�Ћ��A�B�A�B�A�B�A�B�I�J�U���<ډ}ă�;]؉]�������M�3�3�;�~"�U����$    �d$ �t���   ��;�|�U�R�%	  ���E�P�	  ��_^�   [��]Ë��` a a a ��������U��E� �M+]� ���������������U��V��V����`�Hl�AR�Ѓ��Et	V��  ����^]� ���������̡`�H\�������U��`�H\�AV�u�R�Ѓ��    ^]�������������̡`�P\�BQ�Ѓ���������������̡`�P\�BQ�Ѓ����������������U��`�P\�EPQ�J�у�]� ����U��`�P\�EP�EPQ�J�у�]� U��`�P\�EPQ�J�у�]� ���̡`�P\�BQ�Ѓ����������������U��`�P\�EPQ�J �у�]� ����U��`�P\�EP�EPQ�J$�у�]� U��`�P\�EP�EP�EPQ�J(�у�]� ������������U��`�P\�EPQ�J0�у�]� ����U��`�P\�EPQ�J@�у�]� ����U��`�P\�EPQ�JD�у�]� ����U��`�P\�EPQ�JH�у�]� ���̡`�P\�B4Q�Ѓ����������������U��`�P\�EP�EPQ�J8�у�]� U��`�P\�EPQ�J<�у�]� ����U���SVW�}��j �ωu��f�  �`�H\�QV�҃���S���K�  3���~?��I �`�H\�U�R�U��EP�A(VR�ЋM��Q����  �U�R����  ��;�|�_^[��]� �������������U���VW�}�E��P���X�  �}� ��   �`�Q\�BV�Ѓ��M�Q���1�  �E���taS3ۅ�~L�I �UR����  �E�P���
�  �E;E�#���`�Q\P�BV�ЋE����;E��E~߃�;]�|�[_�   ^��]� _�   ^��]� �����������̋�� ����������������������̅�t��j�����̡`�P��  ��`�P��(  ��U��`�P��   ��V�E�P�ҋuP��誨  �M���  ��^��]� ��������̡`�P��$  ��U��`�H��  ]��������������U��`�H���  ]�������������̡`�H��  ��U��`�H���  ]��������������U��`�H��x  ]��������������U��`�H��|  ]��������������U���EV�����t	V��  ����^]� �������������̸   � �������̸   @� �������̸   � �������̸   � ��������U��`�H�QV�uV�҃���^]� �3�� �����������3�� �����������U����   h�   ��@���j P�j �M�Eh�   ��@���R�M��MPQjǅ`���    艺���� ��]���U����   V�u��u3�^��]�h�   ��@���j P�%j �M�U�Eh�   �M���@���Q�U��U��@����ERPj��`���ǅD���k �E���E��o �E�0��E��o �E� �E��o �E�p������� ^��]�������������U���   SV�u(3ۅ��]�u�`�H�A�UR�Ѓ�^3�[��]Ë`�Q�B<W�M3��Ѕ��'  ���  ���E�tq�MQ�M��y�  Wh���M��ˡ��P�M��b�  �u�Wj��U�R�E�P��\���Q�_?腷  ��P��x���R��  ��P�E�P��  ��P����  ���E�t�E� �� t�M����耥  ��t��x�������m�  ��t��\�������Z�  ��t�M̃���J�  ��t�`�Q�J�E�P����у���t�M�� �  �}� t"�U(�E$�M�R�UP�EQ�MRPQ����������U�R��  ����E$�M�UVP�Ej QRP����������`�Q�J�EP�у���_^[��]���������������̋�`����������̋�`����������̋�`�����������U��V�u���t�`�QP��Ѓ��    ^]���������̡`�H��@  hﾭ���Y����������U��E��t�`�QP��@  �Ѓ�]����������������U��`�H���  ]��������������U��`�H��  ]�������������̡`�H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW�qg ������u_^]Ã} tWj V�f ��_������F�d   ^]���U��`�ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW��f ������u_^]�Wj V�f ��_������F�d   ^]�������������U��`�ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW�uf ������u_^]�Wj V�e ��_������F�d   ^]�������������U��`�ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW��e ������u_^]�Wj V�e ��_������F�d   ^]�������������U��`�ɋEt��s�   �I���   j j P�҃�]Ã�s�   VW�xW�ue ������u_^]�Wj V�d ��_������F�d   ^]�������������U��M��t-�=d t�y���A�uP��e ��]á`�P�Q�Ѓ�]��������U��M��t-�=d t�y���A�uP�e ��]á`�P�Q�Ѓ�]��������U��`�H�U�R�Ѓ�]���������U��`�H�U�R�Ѓ�]���������U��`�ɋEt#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�1d ������u_^]�Wj V�Rc ��_������F�d   ^]���������U��`�ɋEtL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]ËMQ������]�������U��E��w�   �`��t�U�IR�URP���   �Ѓ�]Ã�s�   VW�xW�Bc ������u_^]�Wj V�cb ��_������F�d   ^]����������U��E��w�   �`��t,�} �U�IR�URPt���   �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW�b ������u_^]�Wj V��a ��_������F�d   ^]�������U��`�H�U�R�Ѓ�]���������U��`�H�U�R�Ѓ�]���������U��`�H�U�R�Ѓ�]���������U��`�H�U�R�Ѓ�]���������U��`�Hp�]��`�Hp�h   �҃�������������U��V�u���t�`�QpP�B�Ѓ��    ^]���������U��`�Pp�EP�EPQ�J�у�]� U��`�Pp�EP�EPQ�J�у�]� U��`�Pp�EP�EPQ�J�у�]� U��`�Pp�EPQ�J�у�]� ����U���V�u�W�}�����Dz�F�_����D{:�F����$�:b �G��$�]��*b �E���������D{_�   ^��]�_3�^��]���������U��`�P�E���   ��VWP�EP�E�P�ҋu���`�H�QV�ҡ`�H�QVW�ҡ`�H�A�U�R�Ѓ�_��^��]� ������������U���VW�M��0t  �E���}t-�`�Q4P�B�Ѓ����M�u�ht  _3�^��]Ë�R(��`�H0�QW�҃����M�tԋ�R Q�MQ���ҋ�`�P�B �M��Ѓ��t�`�Q0�Jx�E�PW�у��M���s  _��^��]�������U��`�P�B VW�}�����=NIVb��   ��   =TCAbtR=$'  t6=MicM��   �`�Q���   j hIicM���ЋWP�B����_^]� ��BW����_�   ^]� �`�Q���   j hdiem���ЋWP�B����_^]� =INIb��   �~ u���B���F   ��_^]� �~ t���B����_^]� =atniDt5=ckhct=ytsdu?��B����_�F    3�^]� ��B����_^]� 衮��_3�^]� =cnys����_3�^]� ������V�����`�H0�Vh x �҉F���F    ��^�����V��F����t�`�Q0P�B�Ѓ��F    ^�����̡`�P0�A���   P�у����������U��`�P0�E�I���   PQ�҃�]� �������������̡`�I�P0���   Q�Ѓ���������̡`�P0�A���   j j j j j j j j j4P�у�(������̡`�P0�A���   j j j j j j j j j;P�у�(�������U��`�P0�E�IPQ���   �у�]� ��������������U����E V��P�M��q  �`�E�Q�R4Ph8kds�M��ҡ`�E     �H0���   �U R�U�E�P�Ej R�UP�ER�UP�FRj2P�ыu ��(�M���p  ��^��]� ��������������̡`�I�P0���   Q�Ѓ����������U��V��F��u^]� �`�Q0�M ���   j j j j j Q�Mj QjP�ҡ`�H0�U�E���   R�UP�ER�UP�Fj RP�у�D^]� ���̋A��uË`�Q0P�B�Ѓ������̋A��u� �`�Q0P�B�Ѓ�� �U��Q����u�E�    �P��]� �E�H� V�5`�v0Q�MQP���   R�U�R�Ћu�    �F    �`���   j P�BV�Ћ`���   �
�E�P�у�$��^��]� �������U��`�P0�E�I�RPQ�҃�]� �U��A��t)�`�Q0�M���   j j j j j j Qj jP�҃�(]� ���������U��Q��u3�]� �E�H� V�5`�v0Q�MQPR�V�҃�^]� ����������U��Q��u3�]� �E�H� V�5`�v0QP���   R�Ѓ�^]� �����������U��Q��u3�]� �E�H� V�5`�v0Q�MQPR�V\�҃�^]� ����������U��y u3�]� V�u�W�}�؉��ډ�`�P4�A�JhWVP�ы�ډ����ى_^]� �����U��A��u]� �`�Q4�M�RhQ�MQP�҃�]� ����U��A��u]� �`�Q4�M�RpQ�MQP�҃�]� ����U��y u3�]� V�u�W�}�؉��ډ�`�P4�A�JpWVP�ы�ډ����ى_^]� �����U���$VW��htniv�M���l  �`�P�E�R4Phulav�M��ҡ`�P�B4hgnlfhtmrf�M��Ћ`�E�Q�R4Phinim�M��ҡ`�P�E�R4Phixam�M��ҡ`�P�E�R4Phpets�M��ҡ`�P�E�R4Phsirt�M��ҋE =  ��}$u�����t.�`�QP�B4h2nim�M��Ћ`�Q�B4Wh2xam�M��ЋU�M�QR�E�P���K����`���   P�B8�Ћ`���   �
���E�P�у��M���k  _��^��]�  ��������������U���$V��htlfv�M��k  �E�`�P�B,���$hulav�M��Ћ`�E,�Q�R4Phtmrf�M����E�`�P�B,���$hinim�M����E�`�Q�B,���$hixam�M����E$�`�Q�B,���$hpets�M��Ћ`�ED�Q�R4Phsirt�M��������E0��������Dzw���]8����Dzm�؋`�E@�Q�R4Phdauq�M��ҋM�E�PQ�U�R��������`���   P�B8�Ћ`���   �
���E�P�у��M��j  ��^��]�@ �١`�P�B,���$h2nim�M����E8�`�Q�B,���$h2xam�M����V�����U���$V��hgnrs�M���i  �E�`�E��E�   �Q���   �E�Pj�M��ҡ`���   ��U�R�ЋM�`�M����E�   �B���   �M�Qj�M��ҡ`���   ��U�R�ЋU���M�QR�E�P��������`���   P�B8�Ћ`���   �
���E�P�у��M��zi  ��^��]� �U���$V��hCITb�M��i  �`�P�E�R8PhCITb�M��ҡ`�P�E�R4Phsirt�M��ҡ`�P�E�R4Phulav�M��ҋM�E�PQ�U�R�������`���   P�B8�Ћ`���   �
���E�P�у��M���h  ��^��]� U��E��Vj ��P�M�Q�M���  �UPR���)�����`�H�A�U�R�Ѓ���^��]� ����������U��E,��UPj ���T$�$htemf�E$�� �\$�E�\$�E�\$�E�$R�O���]�( �����������U��E,��Pj ���T$�U�$hrgdf�E$�� ����� ������\$�E�����\$�M���\$�E�$R�����]�( ���U��E,��Pj ���T$�U�$htcpf�E$�� �@������\$�E���\$�}�\$�E�$R����]�( ���������������U��Q��u3�]� �E�E�H� V�5`�v0Q�M Q�M���\$�E�$QPR�V(�҃�$^]� ������U��Q��u3�]� �E�H� V�5`�v0Q�MQPR�V,�ҋU3Ƀ�9M^���
]� �������������U��Q��u3�]� �E�H� V�5`�v0Q�MQPR�V,�҃�^]� ����������U��Q��u3�]� �E�H� V�5`�v0Q�MQPR�V0�҃�^]� ����������U��SVW���W��t$�E�H�5`�^0� �uQVP�C0R�Ѓ���u	_^3�[]� �W��t��E�H� �`�[0Q�NQPR�S0�҃���t̋W��tŋE�H� �=`�0Q��VP�G0R�Ѓ���t�_^�   []� ��U��Q��u3�]� �E�H� V�5`�v0Q�MQ�MQPR�V<�҃�^]� ������U��QV3���Wu3��,�E�H� �5`�v0Q�MQPR�V,��3Ƀ�9M������`�M�B�P0VQ�M�ҋ�_^]� ����U��A��Vu3��"�M�Q�	�5`�v0R�URQP�F,�Ѓ����`�Q�E�M�R4PQ�M�ҋ�^]� ���������������U��A����Vu3��"�M�Q�	�5`�v0R�U�RQP�F0�Ѓ����`�E��Q�E�M�R,���$P�ҋ�^��]� �����U�����V���U��V�U����]�Wt$�E�H� �=`�0Q�M�QPR�W0�҃���u
_3�^��]� �V��t�E�H� �=`�0Q�M�QPR�W0�҃���tˋV��tċE�H� �5`�v0Q�M�QPR�V0�҃���t��`�P�M�RH�E�PQ�M��_�   ^��]� �����������U��� ��A���U�V�U��]�Wu3��&�M�Q�	�5`�v0R�U�R�U�RQP�F<�Ѓ����E����}t�`�Q�RH�M�QP���ҋE���t�`�E��Q���$P�B,����_��^��]� U��`�P�E���   Vj ��MP�ҋM$�U Q�MR�Uj Q�MR�UQPR���o���^]�  ����������U��`��P�E���   V���$��MP���E8�E@�M,�Uj P���\$�E0�$Q�E$�� �\$���E�\$�E�\$�$R�K���^]�< ������U��`��P�E���   V���$��MP����Ej j ���T$���$htemf�E$�� �\$�E�\$�E�\$�$P�����^]�$ �����������U��`��P�E���   V���$��MP���E$�Ej �� �\$���E�\$�E�\$�$P�C���^]�$ ��������������U��`��P�E���   V���$��MP����j j ���T$�E�$htcpf�E$�� �@��������\$�E���\$�}�\$�$P����^]�$ ���������������U��`�� V��H�A�U�R�ЋM�E��Qj �U�RP�M�Q�M�����UPR��������`�H�A�U�R�Ћ`�Q�J�E�P�у���^��]� ������������U���dV��M��߆  �`�Q���   P�EP�M�Q�M��P�M��i�  �M�衇  j j �E�P�M��Q�  �MPQ�������`���B�P�M�Q�҃��M��f�  �M��^�  ��^��]� �����U���P��E����]���VW�}��t�`�Q���$P���   �����]���`�U��UЍE��]ȋQ�M���   PQ�E�P���ҋ�M��P�U�H�M�P�U�H�M��P�F���U�u_^��]� �M�E�Q�	�5`�v0R�U R���\$�U��E��$RQP�F(�Ѓ�$_^��]� ���������������U���0�E���M�u�`�H���   �҅�u��]� SVW���k  ��htlfv�MЉu�Z^  �E�}�`�X�U�����$�lK �]��G�$�^K �}�S,�M��$hulav�ҡ`�P�B4hmrffhtmrf�M��Ћ}��`�M�Y���$�K �]��G�$�K �}�S,�M��$hinim�ҋ}��`�M�X���$��J �]��G�$��J �}�S,�M��$hixam����`�P�B,���$hpets�M��Ћ`�Q�B4j hdauq�M��Ћ`�Q�B4Vhspff�M��Ћ`�E �Q�R4Phsirt�M��ҋM�E�PQ�M��U�R�n����`���   P�B8�Ћ`���   �
���E�P�у��M��]  _��^[��]� U��E����V��u�`�H���   �҅�u^��]� ���Ni  �E�F��u3��"�M�Q�	�5`�v0R�U�RQP�F0�Ѓ����E���H��M������\$�M��$��  ��M��P�Q�P�Q�@�A��^��]� ����������U���0��`�]�V���M�]�P���   �E�PQ�M�E�P�ҋ�P�M��Hj �U�P�E P�M��MQ�M�U��UR�U�E�PQR������^��]� ���������������U�����UV�]���E�P�]��ERP�����`�Q�M�R@���E�PQ�M�ҋ�^��]� ����������U��A��u]� �M�Q�	V�5`�v0Rj j j j j j Qj1P���   �Ѓ�(^]� ���������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��A��u]� �`�Q0�M���   j j j j j j j Qj-P�҃�(]� �����U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj j j Q�MQj j j)P�ҋE���(��]� ��U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj j Q�Mj Qj j j)P�ҋE���(��]� ��U��A��u]� �`�Q0�M���   j j j Q�MQ�MQ�Mj Qj/P�҃�(]� ���������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj'P�ҋE���(��]� ������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj,P�ҋE���(��]� ������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�MQ�MQjP�ҋE���(��]� ����������U��`�P0�E�I���   j j j P�EP�EP�Ej Pj.Q�҃�(]� ��������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj:P�ҋE���(��]� ������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj*P�ҋE���(��]� ������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj	P�ҋE���(��]� ��������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj
P�ҋE���(��]� ��������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��A��u]� �`�Q0�M���   j j j Q�MQ�MQ�Mj QjP�҃�(]� ���������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj>P�ҋE���(��]� ������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� �M�Q�	V�5`�v0R�Uj j j j R�URQjP���   �Ѓ�(^]� �����������U����ESVW�M�P�M��(�  �MQ�U�R�M��x�  ��tm�}��E��tN�`���   P�BH�ЋM��I����tQ�W�7�`�[0R�U�j j j j RP���   VjQ�Ѓ�(��t"�MQ�U�R�M���  ��u�_^�   [��]� _^3�[��]� ��������������U��A��u]� �M�Q�	V�5`�v0Rj j j j j j QjP���   �Ѓ�(^]� ���������������U��Q�A��u��]� �`�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� �`�Q0�M�RDQ�MQ�MQP�҃�]� U��A��u]� �`�Q0�M�RHQ�MQ�MQ�MQ�MQ�MQP�҃�]� ���̋A��uË`�Q0P�BX�Ѓ�������U��A��u]� �`�Q0�M�RLQ�MQP�҃�]� ����U��A��u]� �`�Q0�M�RP��   �QP�҃�]� ��U��A��u]� �`�Q0�M�RPQP�҃�]� ��������U��A��u]� �`�Q0�M�RTQ�MQ�MQ�MQP�҃�]� ������������U��`V�u�VW���H4�R�ЋE�F    �~�H� �`�R0Q�MQ���   VP�GP�у�3҅��F_^��]� ���U��A��u]� �`�Q0�M���   j j j j j Qj j jP�҃�(]� �����U��E��u]� �@    �@�I�`�R0P�EPQ���   �у�]� ������̡`�I�P0���   j j j j j j j j j0Q�Ѓ�(�������U��E��u�h� �`�R0�I�R@V�uVP�EPQ�҃�^]� �����������U��`�P0�E�I�RdP�EP�EP�EP�EPQ�҃�]� �U��`�P0�E�I�RpP�EP�EP�EP�EPQ�҃�]� �U��E�P� V�5`�v0R�UR�UR�UR�URP�A�NhP�у�^]� ��������U��E� �`�R0j j j j j j j P�A���   jP�у�(]� �����������U��E� �`�R0j j j j j jj P�A���   jP�у�(]� �����������U��E� �`�R0j j j j j j j P�A���   jP�у�(]� �����������U���V��M��L  �E�H� �`�R0Q�M�Q���   j j j j j P�Fj8P�ы���(��t�M�U�R�L  �M��L  ��^��]� ����������U��E�P� V�5`�v0R�URj j j j j P�A���   j9P�у�(^]� �����U��E�P� V�5`�v0Rj j j j j j P�A���   j"P�у�(^]� �������U��E�P� V�5`�v0Rj j j j j j P�A���   j5P�у�(^]� �������U��E�P� V�5`�v0R�Uj j j j Rj P�A���   j<P�у�(^]� �����U��`�P0�E�I���   j j P�EP�EP�EP�Ej Pj3Q�҃�(]� ������U��`�UVj j j j j R��H0�E�Vj P���   jR�Ћ`�Q0�E�N�RtPQ�҃�0^]� ��U��`�P0�E�I���   j j j j j j Pj jQ�҃�(]� �������������̡`�P0�A���   j j j j j j j j jP�у�(�������U��`�P0�E�I���   j j j j j j j PjQ�҃�(]� �������������̡`�P0�A���   j j j j j j j j j(P�у�(�������U��`�P0�E�I���   j j j j j j P�EPj&Q�҃�(]� ������������U��`�P0�E�I���   j j j j P�EP�Ej Pj+Q�҃�(]� ���������̡`�P0�A���   j j j j j j j j jP�у�(������̡`�P0�A���   j j j j j j j j j#P�у�(�������U��QS�]VW�}���M�t�`�P���   j j���Љ�u��t�`�Q���   j j���Љ�`�Q0�E��H�R`VWQ�҃�_^[��]� �U��`�P0�E�I���   P�EP�EPQ�҃�]� �����̡`�P0�A���   j j j j j j j j j P�у�(������̸   ����������̸   ��������������������������̸   � ��������3�� �����������3���������������� �������������V�����`�H0�Vh x �҉F3��F�F���T��F   ��^�������V��F����t�`�Q0P�B�Ѓ��F    ^������U��E�UVj ��MP�EQ3�9MR��Pj �F    ��
Q��������t�~ t
�   ^]� 3�^]� �U��E�A�I��u3�]� �`�B0Q�H�у�]� ����U��`�P�B S�]V�����=ckhc��   ��   =cksate=TCAb��   �`�Q���   Wj hdiem���Ћ���BSW���F   �Ѓ~ ��t��t��u3Ƀ���Q���C���_^��[]� �~ tK��B����^[]� �~ t6��������t+�F    ^�   []� =atnit�MQS���/���^[]� ^3�[]� �U��V��~ ��   W�}����   �$��� �E;E��   �r�M;M��   �d�U;U��   �V�E;E��   �H�E;E~@;E��   �5�E;E|-;E~v�&�E;E|;E|g��E;E~;E~X��M;MuN�`�M�B0�V���   j j j j j j j QjR���E��(j���\$�E�$W�������F    _^]� Ԧ � � �� � � .� =� L� ����U��V��~ �  �E W�}�E����   �$� � ���]������   �   ���]����A��   �   ���]����A��   �r���]������   �`�E������A��uN��������   �C�E��������u1������A{{�*�E���������E������A�����]����DzU����ء`�U�H0�F���   j j j j j j j RjP���E �U(��(R���\$�E�$W賂�����F    _^]�$ �I �� � $� 6� H� e� ~� �� �� ������������U���E �E�Uj���\$�E�\$�E�$PR�w���]�  ���U���E �E�Uj���\$�E�\$�E�$PR�G���]�  ���U���E �E�Uj���\$�E�\$�E�$PR����]�  ��̋�3�� |��H�H�H�������������VW��3�9~�|�u�`�H4�V�R�Ѓ��~�~_^����U��`�P4�E�I�RtPQ�҃�]� �U��U��t3�A�`�I0R���   P�ҋ`�Q0�M���   QP�҃�]� �`�P0�E�I�R|PQ�҃�]� ������̡`�P4�A�JP�у������������̡`�P4�A�JP�у������������̡`�P4�A�JP�у������������̡`�P4�A�J|P�у������������̡`�P4�A���   P�у����������U��`�P4�E�I�RP�EP�EP�EPQ�҃�]� �����U��`�P4�E�I�RP�EP�EP�EPQ�҃�]� �����U��`�P4�E�I�R PQ�҃�]� �U��`�P4�E�I�R$PQ�҃�]� �U��`�P0�E�I���   P�EP�EP�EPQ�҃�]� ��U��`�P4�E�I���   PQ�҃�]� ��������������U��`�P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U��`�P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U��`�P4�E�I�R(PQ�҃�]� �U��`�P4�E�I�R,P�EP�EPQ�҃�]� ���������U��`�P4�E�I�R0P�EPQ�҃�]� ������������̡`�P4�A�J4P��Y��������������U����UV��EP�M�Q�NR�E�    �E�    �����`�H4�V�AR�Ћ`�Q0�Rhj �M�Q�M�Q�M�Q�M�QP�F�HQ�҃� �} ^t(�} t(�E��M�;�~<�U��;�}3�E�M�;�~)�U���} u�E��M�;�~�U��;�}�   ��]� 3���]� ��������������U��`�P4�E�I�R8PQ�҃�]� �U��`�P4�E�I�R<PQ�҃�]� �U��`�P4�E�I���   P�EPQ�҃�]� ���������̡`�P4�A�J@P�у�������������U��`�P4�E�I�RDP�EPQ�҃�]� �������������U��`�P4�E�I�RHP�EPQ�҃�]� �������������U��`�P4�E�I�RLP�EPQ�҃�]� �������������U��`�P4�E�I�RPP�EPQ�҃�]� �������������U��`SV�uW�����   �QV�҃�����   �`���   �]�QS�҃���SuA�`���   �Q@�ҋء`���   �Q@V�ҋ`�Q4�JPSP�GP�у�_^[]� �`���   �H�у���uD�`���   �H8S�ы`�؋��   �H@V�ы`�J4�WSP�AHR�Ѓ�_^[]� h��h}  ��   �`���   �BV�Ѓ�����   �`���   �]�BS�Ѓ���SuC�`���   �B@�Ћ`���   �؋B8V�Ћ`�Q4�JLSP�GP�у�_^[]� �`���   �H�у���uD�`���   �H8S�ы`�؋��   �H8V�ы`�J4�WSP�ADR�Ѓ�_^[]� h��h�  �
h��h�  �`�Q��0  �Ѓ�_^[]� �U��`�P4�E�I��  P�EP�EP�EPQ�҃�]� ��U��`�P4�E,P�E(P�E$P�E �IP�E�RTP�EP�EP�EP�EP�EPQ�҃�,]�( �������������U��`�P4�E�I�RXP�EP�EP�EPQ�҃�]� ����̡`�P4�A�J`P��Y�������������̡`�P4�A�JdP�у�������������U��`�P4�E�I��   P�EP�EP�EPQ�҃�]� ��U��`�P4�E�I�R\P�EP�EP�EP�EP�EPQ�҃�]� �������������U��`�P4�E�I�RhP�EPQ�҃�]� �������������U��V�u��Wt��؉�}��t��ډ�`�P4�A�JhWVP�у���t��ډ��t��ى_^]� �U��V�u��Wt��؉�}��t��ډ�`�P4�A�JpWVP�у���t��ډ��t��ى_^]� �U��`�P4�E�I�RpP�EPQ�҃�]� �������������U���,V��~ ��   �`�V�H4�AR�Ѓ} t �`�Q0�RlP�F�HQ�҃�^��]� ��hARDb�MԉE��E�    �L8  P�M�Q�N�U�R�����`���   ��U�R�Ѓ��M��]8  ^��]� ������U��`�P4�E�I�RlPQ�҃��   ]� ������������U��`�E�P4�E�I���   P�E���\$�E�$PQ�҃�]� ����������U��`�P4�E�I���   P�EP�EPQ�҃�]� �����̡`�P4�A���   P�у���������̸   ����������̸   �����������U��`V��H4�V�A$h�  R�Ћ`�Q4�E�MP�EQ�MP�FQ�JP�у�2�^]� ��������U��U��@R�UR�UR�UR��]� �̸   � ��������3�� ������������ �������������3�� ������������ �������������U��`�P4�E�I�RxP�EP�EP�EPQ�҃�]� �����U��`�P0�E�I�I���   P�EP�EPQ�҃�]� ���U��QS�]VW�}���M�t�`�P���   j j���Љ�u��t�`�Q���   j j���Љ�`�Q4�E��H�RpVWQ�҃�_^[��]� �U��Q�`�P�B SVW�}���3���=INIb�/  �  =SACbvt+=$'  t
=MicM�  ��B$W����_�   ^��[��]� ��R3��E��E�EP�M�Q���҅�t�`�U�H4�E�R�VP�AR�Ѓ�_�   ^��[��]� =ARDb�  �`�Q���   j j���Ћ`�Qj �؋��   j���Ћ`�Qj �E����   j���Ћ`�Qj �E���   j���ЋM���RWP�EPQS����_�   ^��[��]� ��P����_�   ^��[��]� =NIVbetJ=NPIbt0=ISIbu\�>���Y���P���1���P�G����_�   ^��[��]� ��BW����_^[��]� ��B����_�   ^��[��]� =cnyst_^��[��]� �`�Q���   j hIicM���ЋWP�B ����_^[��]� �������������U��`�P4�E�I�RTh����h����h����P�EP�Eh����h����h����h����PQ�҃�,]� ������U���V��hYALf�M��*3  �`�Q4�JlP�FP�у��M��L3  ^��]��������V�����`�H0�Vh x �҉F���F    ���F   ��^��������V��F����t�`�Q0P�B�Ѓ��F    ^������U��`�P�B VW�}�����=cksat`=ckhct�MQW��譾��_^]� �Nj j j j j j �F   �`�B0���   j j j Q�҃�(��t'_�F    �   ^]� �~ t��P����_^]� _3�^]� ���U��`�H���  ]��������������U��`�H0���   ]��������������U��`�H0�U�E��VWRP���   �U�R�Ћ`�Q�u���BV�Ћ`�Q�BVW�Ћ`�Q�J�E�P�у�_��^��]������������U��`�H0���   ]��������������U��`�H0���   ]��������������U��Ej0P�k����]��������������U��Ej0P�r!  ��P��j����]�����U��E�M��j0PQ�U�R�w!  ��P�j���`�H�A�U�R�Ѓ���]�������U��E�M�U��j0PQR�E�P�"  ��P�zj���`�Q�J�E�P�у���]��U��Ej$P�Rj��3Ƀ�������]����U��Ej$P�   ��P�)j��3Ƀ�������]�����������U��E�M��Vj$PQ�U�R�   ��P��i���`3Ƀ��B�P����M�Q�҃���^��]��������U��E�M�U��Vj$PQR�E�P��!  ��P�i���`3Ƀ��B�P����M�Q�҃���^��]����U��`�H�U�E���   RPj �у�]���������������U��`�H�U�ER�UP���   Rj �Ѓ�]�����������U��`�P4�E�I�R,P�EP�EPQ�҃�]� ���������U��`�P4�E�I�R0P�EPQ�҃�]� ������������̡`�P4�A�J4P��Y��������������U��U��V��EP�M�QR���d����`�H0�E�P� R�U�R�U�R�U�R�U�R�VP�AhR�Ѓ��} ^t(�} t(�E�M�;�~<�U��;�}3�E�M�;�~)�U���} u�E�M�;�~�U��;�}�   ��]� 3���]� �����������U��E��SVW��u�Y�`�P�}���   j hdiuM���Ћ���tK;3u	_^3�[]� �`�Q���   j hIicM����;�u�`�Q���   j h1icM���Шu��3_^�   []� �����U��`�P�BT��(V�uhfnic���Ѕ�t�`�Q�ȋ��   j
�Ѕ���   �`�Q�RPhfnic�E�P����P�M���,  �M��-  �u�E�P���	-  �M���,  �`�Q�B ���Ѓ��t�`�Q�B ���Ѕ�u�`�Q�B$hfnic���Ћ`�E�Q�R8Pj
����^��]���������U��`�P0�E�IP�EP�EP�EPQ���   �у�]� ��U��`�P0�E�IV�p� ���   V�uj j j V�uVj Pj=Q�҃�(^]� ����U��`�P0�E�IV�p� ���   V�uV�uj j j�Vj Pj=Q�҃�(^]� ���̡`�I�P0���   j j j j j j j j j6Q�Ѓ�(�������U��V�����`�H0�WVh x �ҋ}�F�E�F    �F   ���F�`�Q���   ��j hmyal���Ѓ��Ft��t�F    �`�Q���   j
hhfed���ЉF_��^]� �����������U��`�P�B VW�}�����=ytsdt�MQW������_^]� �`�B0�N���   Q�ҋ�P������_�   ^]� ��3���������������3�������������������������������3���������������3���������������3���������������3�� �����������U��V���PD�҅�t�E9Ft�F��PH����^]� �����̋A������������̋A��uË ��������������������̸h������������U���E�Y(]� ���U���(V���P(�M�Q���ҋN��t&�`�R0j j j j j j P���   j jQ�Ѓ�(�`�Q�J�E�P�ы`�B�P�M�Q�ҋF����t �`�Q0�RHj �M�Qj jj?j P�҃��`�H�A�U�WR�Ћ`�Q�J�E�P�ыF����u3��;�`�E�    �J0�U�Rj j j h  
 j�U�Rh�  jP���   �Ћ}���(�`�Q�J�E�P�у���_u3�^��]Ë`�B�P�M�Q�ҋF����t �`�Q0�RHj �M�Qj j j8j P�҃��`�H�A�U�R�ЋF����t�`�Q0jP�BP�Ѓ��`�Q�J�E�P�у��M��'  Ph   h  K j;�U�Rh	��h�  ��跶���`�H�A�U�R�Ѓ��M���'  �F��t�`�Q0P�BX�Ѓ��F��t�`�Q0P�BX�Ѓ��F��t'�`�Q0j j j j j jj j jP���   �Ѓ�(j�v$��`�����   ^��]�����U���SV��W�~j���y�  ��V�^(3ۉ^4�^8�^<�`�H0�Ah�   R�Ћ`�Q�J�E�P�ы`�B�PSj��M�hx�Q�҃�SS�E�P�M�Q���E��  �]��i����`�B�P�M�Q�҃�Sj��躱  _^[��]���̍A�������������U��VW��~4 tA�I �`�H��0  h��hj  ��j
��i���`�HP�V �AR�Ѓ���uQ9F4u`�QP�Bh�~0���Ѓ~4 t;�`�Q��0  h��h�  �Ћ`�QP�Bl�������m���_3�^]� �M�U�N8�V4�`�PP�Bl�~0���Ѓ~4 t%j
�3i���`�QP�F �JP�у���u�9F4uۋ`�BP�PhS���ҋ^<�F<    �`�PP�Bl���Ћ�[_^]� ��U��`�P�B ��@VW�}�����=MicMtI=fnic��   j�M��%  �uP���M%  �M��5%  �`�Q�B4jj����_�   ^��]� �`�Q���   j hIicM����=�����   htats�M��$  �`�Q�B0j j�M��ЍM�Q�U�R�E�P���E��  �E�    �̴���`���   �
�E�P�у��M��$  �F���F   t�`�J0�QP�҃��EPW���a���_^��]� ���������U��E��V��t3�^]� j�N�a�  j�]���F    �v����t�`�H0�QV�҃��   ^]� ��������������j����  j�_]����3�����������U��E3�h�����h  ���P�Ej ��R�Uj PR�s���]� ���������������U��Q�Q��u3���]� �E�H� V�5`Q�M�Q�E�    �v0PR�V8�ҋ�����t@�E���t9�`�Q�M�RQP�ҋE�����t�`�QW��P�B��W�s�����_��^��]� ������U��`��V��H�A�U�R�ЋU���M�QR���D�������u�`�H�A�U�R�Ѓ�3�^��]� �M�Q�M�UK  �`�B�P�M�Q�҃���^��]� �������U��`��V��H�A�U�R�ЋU���M�QR��������M��`�P�R8�E�PQ�M�ҡ`�H�A�U�R�Ѓ���^��]� �������������U���V��M��H  �M�E�PQ��������`���B�U�@<�M�Q�MR�ЍM��]I  ��^��]� ����U��`�P�E���   Vj ��MP��h���h  �j j jj P�EP���S���^]� ��������������U��`V�uW�����   �QV�҃���Vu,�`���   �Q@�ҋ`�Q4�J P�GP�у�_^]� �`���   �H�у���u.�`���   �H8V�ы`�J4�WP�A$R�Ѓ�_^]� �`�Q��0  h��h	  �Ѓ�_^]� �����U���4�`�H�QSVW�}W�ҡ`�P�u���   ��3�SS�Ή]�Ћ`�QS�E����   j���Ћ�;��M  �d$ �} ~l�`�Q�J�E�P�ы`�B�Pj j��M�h|�Q�ҡ`�P�B<�����Ћ`�Q�RLj�j��M�QP���ҡ`�H�A�U�R�Ѓ��`�Q0�E����   VP�M�Q�ҋ�`�H�A�U�R�Ћ`�Q�J�E�PV�ы`�B�P�M�Q�ҡ`�P�B<�����Ћ`�Q�RLj�j��M�QP���ҡ`�H�A�U�R�Ћ`�Q�u���   �E��j ��
S���Ћ`�Q���   �E�j �CP���ҋ����������_^[��]���������������U��E�PV��3Ƀ8������t�   3�h�����h  ���Pj ��Qj R�UR���{���^]� ������U��E3҃8�@V�u ��V�uVR�UR�UR�UR�UPR�?���^]� ����������U��E�E43҃8��R�U<R�U(���\$�E,�$R�E �� �\$�E�\$�E�\$�@�E�$P�2���]�8 ��������������U��E�@3҃8��E��Rj ���T$�$htemf�E �� �\$�E�\$�E�\$�$P�ױ��]�  ���U��E�E 3҃8��R�� �\$�E�\$�E�\$�@�E�$P�Z���]�  ������U��E�@3҃8��E��Rj ���T$�$htcpf�E �� �@������\$�E���\$�}�\$�$P�;���]�  �������U��E3҃8��R�UR�UR�UR�UP�EPR����]� U��E3҃8V�u��V��RP�EP�O���^]� ����������U��Q��u3�]� �E�E�H� V�5`�v0Q�M Q�M���\$���E�$QPR�V(�҃�$^]� ���U��`�P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U��`�P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U��`��P�E���   V���$��MP�ҋ���u�^�    ^]� ��u�^����D{�   ^]� ��^]� ������U���0��`�U�V�U���M�]�P���   �E�PQ�M�E�P�ҋ���̉�P�Q�P�Q�P�Q�P�@�Q�A����  ^��]� ��������U��� ��`�]�V���M�]��P���   �E�PQ�M�E�P�ҋ���̉�P�Q�P�@�Q�A����  ^��]� �����U���VW�};}�M�us�`�P�u���   j htsem���Ѕ�uS�`�QP���   hrdem���Ѕ�u6�MQ�M�U�R�E�}�E�������t�E�M�P�w  _�   ^��]� _3�^��]� U���VW�};}�M�us�`�P�u���   j htsem���Ѕ�uS�`�QP���   hrdem���Ѕ�u6�MQ�M�U�R�E�}�E��ײ����t�E�M�P��  _�   ^��]� _3�^��]� U���SVW�};}��uz�`�P�u���   j htsem���Ѕ�uZ�`�QP���   hrdem���Ѕ�u=��M�Q�]��M�U�R�}��E�腲����t�E������$�  _^�   [��]� _^3�[��]� ��������U���4�ESW�};ǉM�t;Et	;E��   �`�P�]���   j htsem���Ѕ���   �`�QP���   hrdem���Ѕ�uj�M��U�U܉E��UԉE��]̉E�M�E�P�M�Q�M�U�U�R�E�P�}�������t+�E̋M�������E��X�E��X��  �   _[��]� _3�[��]� ��������U���SVW�};}����   �`�P�u���   j htsem���Ѕ�uj�`�QP���   hrdem���Ѕ�uM��U�M��]���Q�M�]��E�R�E�P�}��h�����t%�E��������E��X�  �   _^[��]� _^3�[��]� ���̋A���X(Q�ȋB$��j j h����pS�����������������U��`��0VW���H�A�U�R�Ћ`�Q�J�E�P�ыE���U�RP�M�Q�M輡���`�J�U�RP�A�Ћ`�Q�J�E�P�ы`�B�P�M�Q�ҡ`�H�Q��V�ҡ`�H�A�U�VR�Ѓ�����  �`�Q�J�E�P�у�_^��]� ������������U���SVW�};}����   �`�P�u���   j htsem���Ѕ�ue�`�QP���   hrdem���Ѕ�uH�`�Q�J�E�P�ыM���U�R�E�P�}��E�    �-�����u �`�Q�J�E�P�у�3�_^[��]� ���U��R��8�����  �`�H�A�U�R�Ѓ�_^�   [��]� ��U��V�u���  ��^]� �����������U���L�`SV��H�A�U�R�Ћ`�Q�J3�Sj��E�h��P���F(�@���S�U�SR�E��  �]��h�  P�E�P�8����P�M�Q�J����P�U�R���R����`�H�A�U�R�Ћ`�Q�J�E�P�ы`�B�P�M�Q�҃�htats�M��=  �`�P�B0jj�M����F(�`�Q�B,���$j�M��ЍM�Q�U�R�E�P���E��  �]��P����`���   �
�E�P�у�9^4t^�`�BP�PhW�~0���ҋF4;�t�N8Q�Ѓ��F<�^8�^4��`�B��0  h��h�  �у��`�BP�Pl����_�M��  ^[��]� ������U�����u�E�    �A]� ��u�Q;Ut�   ]� U�����u�E�    �Y]� ��u�E�Y����D{�   ]� �����������U�����u�E�    �Y�E�Y�E�Y]� ��u-�E�Y����Dz�E�Y����Dz�E�Y����D{�   ]� �����U��V�����u#�E�M�U�F�E�N�V�    �F^]� ��u�MQ�VR��������t�   ^]� �������������U��V��~ �|�u�`�H4�V�R�Ѓ��E�F    �F    t	V葘������^]� �������U��V��F����t�`�Q0P�B�Ѓ��E�F    t	V�H�������^]� ��������������U���V��3ɍF��H������`�M��M����   �RQ�M�QP�ҡ`���   ��U�R�Ѓ���^��]��������������U��V�����u �    �`�H�A���UVR�Ѓ��#��u�`�Q�Rx�EP�N�҅�t�   �`�H�A�UR�Ѓ�^]� �������U��E��u�h�MP�EPQ��  ��]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3h��j;h�j轗������t
W����7  �3����Fu_^]� �~ t3�9_��^]� �`�H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   �`�H<�Q��3Ʌ����^��������������̃y t�   ËA��uË`�R<P��JP�у��������U����u�`�H�]� �`�J<�URP�A�Ѓ�]� ���������������U��h��u�`�H�]Ë`�J<�URP�A�Ѓ�]�U��h��$��Vu�`�H�1��`�J<�URP�A�Ѓ����`�Q�J�E�SP�ы`�B�P�M�QV�ҡ`�H�A�U�R�Ћ`�Q�Jj j��E�h̵P�ы`�B�@@�� j �M�Q�U�R�M��Ћ`�Q�J���E�P���у���[t.�`�B�u�HV�ы`�B�P�M�Q�҃���^��]á`�P�E��RHjP�M��ҡ`�P�E�M��RLj�j�PQ�M��ҡ`�H�u�QV�ҡ`�H�A�U�VR�Ћ`�Q�J�E�P�у���^��]���������������U��h��$��SVu�`�H�1��`�J<�URP�A�Ѓ����`�Q�J�E�P�ы`�B�P�M�QV�ҡ`�H�A�U�R�Ћ`�Q�Jj j��E�h̵P�ы`�B�@@�� j �M�Q�U�R�M��Ћ`�Q�J���E�P���у���t/�`�B�u�HV�ы`�B�P�M�Q�҃���^[��]á`�P�E��RHjP�M��ҡ`�P�E�M��RLj�j�PQ�M��ҡ`�H�A�U�R�Ћ`�Q�Jj j��E�h̵P�ы`�B�@@��j �M�Q�U�R�M��Ћ`�Q�J���E�P���у����3����`�P�E��RHjP�M��ҡ`�P�E�M��RLj�j�PQ�M��ҡ`�H�u�QV�ҡ`�H�A�U�VR�Ћ`�Q�J�E�P�у���^[��]����������������U��h��$��SVu�`�H�1��`�J<�URP�A�Ѓ����`�Q�J�E�P�ы`�B�P�M�QV�ҡ`�H�A�U�R�Ћ`�Q�Jj j��E�h̵P�ы`�B�@@�� j �M�Q�U�R�M��Ћ`�Q�J���E�P���у���t/�`�B�u�HV�ы`�B�P�M�Q�҃���^[��]á`�P�E��RHjP�M��ҡ`�P�E�M��RLj�j�PQ�M��ҡ`�H�A�U�R�Ћ`�Q�Jj j��E�h̵P�ы`�B�@@��j �M�Q�U�R�M��Ћ`�Q�J���E�P���у����3����`�P�E��RHjP�M��ҡ`�P�E�M��RLj�j�PQ�M��ҡ`�H�A�U�R�Ћ`�Q�Jj j��E�h̵P�ы`�B�@@��j �M�Q�U�R�M��Ћ`�Q�J���E�P���у���������`�P�E��RHjP�M��ҡ`�P�E�M��RLj�j�PQ�M��ҋu�E�P����,���`�Q�J�E�P�у���^[��]�������U��h��$��SVu�`�H�1��`�J<�URP�A�Ѓ����`�Q�J�E�P�ы`�B�P�M�QV�ҡ`�H�A�U�R�Ћ`�Q�Jj j��E�h̵P�ы`�B�@@�� j �M�Q�U�R�M��Ћ`�Q�J���E�P���у���t/�`�B�u�HV�ы`�B�P�M�Q�҃���^[��]á`�P�E��RHjP�M��ҡ`�P�E�M��RLj�j�PQ�M��ҡ`�H�A�U�R�Ћ`�Q�Jj j��E�h̵P�ы`�B�@@��j �M�Q�U�R�M��Ћ`�Q�J���E�P���у����3����`�P�E��RHjP�M��ҡ`�P�E�M��RLj�j�PQ�M��ҡ`�H�A�U�R�Ћ`�Q�Jj j��E�h̵P�ы`�B�@@��j �M�Q�U�R�M��Ћ`�Q�J���E�P���у���������`�P�E��RHjP�M��ҡ`�P�E�M��RLj�j�PQ�M���j h̵�M��b*���`�P�R@j �E�P�M�Q�M��҅��`�H�A�U�R���Ѓ���t/�`�Q�u�BV�Ћ`�Q�J�E�P�у���^[��]Ë`�M��B�PHjQ�M��ҡ`�P�E�M��RLj�j�PQ�M��ҋu�E�P���)���`�Q�J�E�P�у���^[��]���������������U��`�H<�A]����������������̡`�H<�Q�����V��~ u>���t�`�Q<P�B�Ѓ��    W�~��t���J-  W�������F    _^��������U���V�E�P����>  ��P��������M���	-  ��^��]��̃=p uK�h��t�`�Q<P�B�Ѓ��h    �t��tV����,  V芋�����t    ^������������U���8�`�H�AS�U�V3�R�]��Ћ`�Q�JSj��E�hеP�ы`�B<�P�M�Q�ҋ�`�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��h�  �M�Q�U�R�M�踎  ����   W�}�}���   �`���   �U��ATR�Ћ�����tB�`�Q�J�E�P���у��U�Rj�E�P�������`�Q�ȋBxW�Ѕ��E�t�E� ��t�`�Q�J�E�P����у���t�`�B�P�M�Q����҃��}� u"�E�P�M�Q�M���  ���;����E�_^[��]ËU��U�_�E�^[��]��������������U���DSV�u3�;�]�u_�`�H�A�U�R�Ћ`�Q�JSj��E�hеP�ы`�B<�P�M�Q�ҋ�`�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]���  �M�Q�U�R�M��1�  ���p  W�}��I �E����   �`���   �U��ATR�Ћ�������   �`�Q�J�E�P���ы`�B���   ���M�Qj�U�R���Ћ`�Q�J���E�P�ы`�B�P�M�QV�ҡ`�H�A�U�R�Ћ`�Q�Bx��W�M��Ѕ��Et�E ��t�`�Q�J�E�P����у���t�`�B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*�`���   P�BH�Ћ`�Q���ȋBxW�Ѕ�t"�M�Q�U�R�M��ҋ  ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M��3�  �EP�M�Q�M�u��u�}�  ����   �u���E���tA��t<��uZ�`���   �M�PHQ�ҋ`�Q���ȋBxV�Ѕ�u-�   ^��]Ë`���   �E�JTP��VP�[�������uӍUR�E�P�M���  ��u�3�^��]����������V��~ u>���t�`�Q<P�B�Ѓ��    W�~��t���
(  W�Ԇ�����F    _^�������̡`�P�BVj j����Ћ�^���������U��`�P�E�RVj P���ҋ�^]� U��`�P�E�RVPj����ҋ�^]� �`�P�B�����U��`�P���   Vj ��Mj V�Ћ�^]� �����������U��`�P�EPQ�J�у�]� ����U��`�P�EPQ�J�у������]� �������������U��`�P�E�RtP�ҋ`���   P�BX�Ѓ�]� ���U��`�P�E�Rlh#  P�EP��]� ���������������U��`�P�E�RlhF  P�EP��]� ���������������U��`�P�E�RtP�ҋ`���   �M�R`QP�҃�]� ���������������U��`�P���   ]��������������U��`�P�E���   P�҅�u]� �`���   P�B�Ѓ�]� �������̡`�HL���   ��U��`�H@�AV�u�R�Ѓ��    ^]�������������̡`�HL�������U��`�H@�AV�u�R�Ѓ��    ^]�������������̡`�PL���   Q�Ѓ�������������U��`�PL�EP�EPQ���   �у�]� �������������U��`V��HL���   V�҃���u�`�U�HL���   j RV�Ѓ�^]� �`���   �ȋBP�Ћ`���   �MP�BH��^]� �����̡`�PL��(  Q�Ѓ�������������U��`�PL�EP�EPQ��,  �у�]� ������������̡`�HL�Q�����U��`�H@�AV�u�R�Ѓ��    ^]��������������U��`�PL�E�R��VPQ�M�Q�ҋu��P���%����M��=�����^��]� ����U��`�PL�EPQ���   �у�]� �U��`�PL�EP�EPQ�J�у�]� �`�PL�BQ�Ѓ���������������̡`�PL�BQ�Ѓ���������������̡`�PL�BQ�Ѓ����������������U��`�PL�EP�EP�EPQ�J �у�]� ������������U��`�PL�EPQ��4  �у�]� �U��`�PL�EP�EP�EPQ�J$�у�]� ������������U��`�PL�EP�EP�EP�EPQ�J(�у�]� �������̡`�PL�B,Q�Ѓ���������������̡`�PL�B0Q�Ѓ����������������U��`�PL�EP�EPQ��  �у�]� ������������̡`�PL���   Q�Ѓ�������������U��`�PL�E��  ��VPQ�M�Q�ҋu��P�������M�������^��]� ̡`�PL�B4Q�Ѓ���������������̡`�PL�B8j Q�Ѓ��������������U��`�PL���   ]��������������U��`�PL���   ]��������������U��`�PL���   ]��������������U��`�PL���   ]��������������U��`�PL���   ]��������������U��`�PL���   ]��������������U��`�PL���   ]��������������U��`�PL���   ]��������������U��`�PL���   ]��������������U��`�PL�EPQ�J<�у�]� ���̡`�PL�BQ��Y�U��`�PL�EP�EPQ�J@�у�]� U��`�PL�Ej PQ�JD�у�]� ��U��`�PL�Ej PQ�JH�у�]� ��U��`�PL�EjPQ�JD�у�]� ��U��`�PL�EjPQ�JH�у�]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}�贔  W�M�Q�U�R��褛  ���M�����  ��t�`���   ��U�R�Ѓ�_^3�[��]Ë`���   �J8�E�P�ы`�����   ��M�Q�҃�_��^[��]��������������U���$3�V�E��E�E��P�M��E�   �E�   �E��  ���  j�M�Q�U�R����  �M��e�  �`���   ��U�R�Ѓ�^��]�����������U���$�`�UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��z�  j�E�P�M�Q��艚  �M���  �`���   ��M�Q�҃�_^��]� ��U���$�`�UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}����  j�E�P�M�Q���	�  �M��a�  �`���   ��M�Q�҃�_^��]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}�蔒  W�M�Q�U�R��脙  ���M������  ��t+�u���	  �`���   ��U�R�Ѓ�_��^[��]� �`���   �JL�E�P�ыu��P���u  �`���   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��ԑ  W�M�Q�U�R���Ę  ���M����7�  ��t+�u���I  �`���   ��U�R�Ѓ�_��^[��]� �`���   �JL�E�P�ыu��P���  �`���   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}���  W�M�Q�U�R����  ���M����w�  _^��[t�`���   ��U�R�������]Ë`���   �J<�E�P���]��`���   ��M�Q���E�����]���������������U���$SVW3��E��P�M��}܉}��E��  �}��}��d�  W�M�Q�U�R���T�  ���M����ǂ  ��t�`���   ��U�R�Ѓ�_^3�[��]Ë`���   �J8�E�P�ы`�����   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}�贏  W�M�Q�U�R��褖  ���M�����  ��t-��u�`����   ���^�U�R�Ѓ�_��^[��]� �`���   �JP�E�P�ы�u�H��P�@�N�`�V���   �
�F�E�P�у�_��^[��]� �����̡`�PL���   Q��Y��������������U��`�PL�E���   ��jPQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U��`�PL�E���   ��j PQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���$SVW3��E��P�M��}܉}��E��  �}��}��$�  W�M�Q�U�R����  ���M���臀  ��t-��u�`����   ���^�U�R�Ѓ�_��^[��]� �`���   �JP�E�P�ы�u�H��P�@�N�`�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��T�  W�M�Q�U�R���D�  ���M����  ��t-��u�`����   ���^�U�R�Ѓ�_��^[��]� �`���   �JP�E�P�ы�u�H��P�@�N�`�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}�脌  W�M�Q�U�R���t�  ���M�����~  ��t-��u�`����   ���^�U�R�Ѓ�_��^[��]� �`���   �JP�E�P�ы�u�H��P�@�N�`�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}�贋  W�M�Q�U�R��褒  ���M����~  ��t�`���   ��U�R�Ѓ�_^3�[��]Ë`���   �J8�E�P�ы`�����   ��M�Q�҃�_��^[��]��������������U����E3�V�]�E��E��E��P�M�E�   �E��  ���  j�M�Q�UR����  �M�f}  �`���   ��U�R�Ѓ�^��]� ���������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E�菊  j�U�R�E�P��螑  �M���|  �`���   �
�E�P�у�^��]� ��������U���$�`�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��
�  j�E�P�M�Q����  �M��q|  �`���   ��M�Q�҃�_^��]� ��U���$�`�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}�芉  j�E�P�M�Q��虐  �M���{  �`���   ��M�Q�҃�_^��]� ��U���$�`�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��
�  j�E�P�M�Q����  �M��q{  �`���   ��M�Q�҃�_^��]� ��U���$�`�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}�芈  j�E�P�M�Q��虏  �M���z  �`���   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E���  j�U�R�E�P���.�  �M��z  �`���   �
�E�P�у�^��]� ��������U���$SVW3��E��P�M��}܉}��E��  �}��}�贇  W�M�Q�U�R��褎  ���M����z  ��t-��u�`����   ���^�U�R�Ѓ�_��^[��]� �`���   �JP�E�P�ы�u�H��P�@�N�`�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}���  W�M�Q�U�R���ԍ  ���M����Gy  ��t�`���   ��U�R�Ѓ�_^3�[��]Ë`���   �J8�E�P�ы`�����   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��4�  W�M�Q�U�R���$�  ���M����x  ��t�`���   ��U�R�Ѓ�_^3�[��]Ë`���   �J8�E�P�ы`�����   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ����U���$�`�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��J�  j�E�P�M�Q���Y�  �M��w  �`���   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��߄  j�U�R�E�P����  �M��Fw  �`���   �
�E�P�у�^��]� ��������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��o�  j�U�R�E�P���~�  �M���v  �`���   �
�E�P�у�^��]� ��������U��`�H���   ]��������������U��`�H���   ]�������������̡`�H���   ��`�H���   ��U��`�H���   V�u�R�Ѓ��    ^]�����������U��`�H���   ]��������������U��`�HL�QV�ҋ���u^]á`�H�U�ER�UP���  RV�Ѓ���u�`�Q@�BV�Ѓ�3���^]����������U��`�H�U�E���  R�U�� P�ERP�у�]������U��`�H���   ]��������������U��`�H�U �ER�UP�ER�UP�ER�UP���   R�Ѓ�]������������̡`�PL�BLQ�Ѓ���������������̡`�PL�BPQ�Ѓ����������������U��`�PL�EP�EPQ�JT�у�]� U��`�PL�EPQ��  �у�]� �U��`�PL�EPQ���   �у�]� ̡`�PL�BXQ�Ѓ����������������U��`�PL�EP�EP�EPQ�J\�у�]� ������������U���4�`SV��HL�QW�ҋ�3�;��}��x  �M������`�E�EԋE�]Љ]؉]܉]�]��}̋Q�R0Ph]  �M��ҡ`���   �BSSW���Ѕ���   �`�QL�BW�Ћ���;���   ��    �`���   �B(���ЍM�Qh�   ���u�� ��������   �M�;���   �`���   ���   S��;�tm�`���   �ȋB<V�Ћ`���   ���   �E�P�у�;�t�`�B@�HV�у�;����\����}��M��4���M��I�����_^[��]� �}��`�B@�HW�ы`���   ���   �M�Q�҃��M��94���M�����_^3�[��]� �����̡`�PL�B`Q�Ѓ���������������̡`�PL�BdQ�Ѓ����������������U��`�PL�EPQ�Jh�у�]� ���̡`�PL��D  Q�Ѓ������������̡`�PL�BlQ�Ѓ����������������U��`�PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U$�EV�Eh�
h�
h�
h�
R�Q�U R�UR�UR�U���A�$�5`�vLRP���   Q�Ѓ�4^]�  ������̡`�PL���   Q�Ѓ�������������U��`�PL�EP�EP�EPQ��   �у�]� ���������U��`�PL��H  ]�������������̡`�PL��L  ��U��`�PL��P  ]��������������U��`�PL��T  ]��������������U��`�PL�EP�EP�EP�EP�EPQ���   �у�]� �U��`�PL�EP�EP�EPQ���   �у�]� ���������U��`�PL�EP�EP�EP�EPQ��   �у�]� �����U��`�HL���   ]��������������U��`�HL���   ]��������������U��`�HL���   ]�������������̡`�HL��  ��`�HL��@  ��h�Ph^� ���  ���������������U��Vh�j\h^� ��蹇  ����t�@\��t
�MQV�Ѓ�^]� ������������U��� �`V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ};��E�t`;�t\�`�QLjP���   ���ЋM��U�Rh=���M�}�������`���   ���   �U�R�Ѓ��M��u���/����_^��]Ë`���   ���   �E�P�у��M��u��/��_�   ^��]����U��� �`V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ};��E�t`;�t\�`�QLjP���   ���ЋM��U�Rh<���M�}��������`���   ���   �U�R�Ѓ��M��u���.����_^��]Ë`���   ���   �E�P�у��M��u���.��_�   ^��]���̡`V�񋈈   ���   V�҃��    ^��������������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������U���   V���P  �����   �ESP�M��H  �`�Q�J�E�P�ы`�B�Pj j��M�h��Q�҃��E�P�M��  j j��M�Q�U�R��d���P�4  ��P�M�Q��  ��P�U�R�  ���P�Q  ���M����A  �M��9  ��d����.  �M��&  �`�H�A�U�R�Ѓ��M��
  ��[t	V��O  ����^��]� ���U��EVP���QY  �����^]� �����Q�O  Y���������U��E�M�U�H4�M�P �U��M�@k �@8��@<p��@@�o �@D�o �@H �@L0��@P��@l@��@X �@\��@`�@d��@T�o �@h���@p��@t��P0�H(�@,    ]��������������U���   h�   ��`���j P�4�  �M�U�Ej Q�MRPQ��`���R�����E �Uh�   ��`���Q�E��ERPj�%����8��]��������������̋�`<����������̋�` ����������̋�`@����������̋�`����������̋�`4����������̋�`����������̋�`8����������̋�`,�����������U��`�P�EP�EP�EPQ�J�у�]� �����������̡`V��H�QV�ҡ`�H$�QDV�҃���^�����������U��`V��H�QV�ҡ`�H$�QDV�ҡ`�U�H$�AdRV�Ѓ���^]� ��U��`V��H�QV�ҡ`�H$�QDV�ҡ`�U�H$�ARV�Ѓ���^]� ��U��`V��H�QV�ҡ`�H$�QDV�ҡ`�H$�U�ALVR�Ѓ���^]� �̡`V��H$�QHV�ҡ`�H�QV�҃�^�������������U��`�P$�EPQ�JL�у�]� ����U��`�P$�R]�����������������U��`�P$�Rl]����������������̡`�P$�Bp����̡`�P$�BQ�Ѓ����������������U��`�P$��VWQ�J�E�P�ы`�u���B�HV�ы`�B�HVW�ы`�B�P�M�Q�҃�_��^��]� ���U��`�P$�EPQ�J�у�]� ����U��`�P$��VWQ�J �E�P�ы`�u���B�HV�ы`�B$�HDV�ы`�B$�HLVW�ы`�B$�PH�M�Q�ҡ`�H�A�U�R�Ѓ� _��^��]� ���U��`�P$��VWQ�J$�E�P�ы`�u���B�HV�ы`�B$�HDV�ы`�B$�HLVW�ы`�B$�PH�M�Q�ҡ`�H�A�U�R�Ѓ� _��^��]� ���U���V�uV�E�P�l������e����`�Q$�JH�E�P�ы`�B�P�M�Q�҃���^��]� ����̡`�P$�B(Q��Yá`�P$�BhQ��Y�U��`�P$�EPQ�J,�у�]� ����U��`�P$�EPQ�J0�у�]� ����U��`�P$�EPQ�J4�у�]� ����U��`�P$�EPQ�J8�у�]� ����U��`�UV��H$�ALVR�Ѓ���^]� ��������������U��`�H�QV�uV�ҡ`�H$�QDV�ҡ`�H$�U�ALVR�Ћ`�E�Q$�J@PV�у���^]�U��`�UV��H$�A@RV�Ѓ���^]� ��������������U��`�P$�EPQ�J<�у�]� ����U��`�P$�EPQ�J<�у������]� �������������U��`�P$�EP�EPQ�JP�у�]� U��`�P$�EPQ�JT�у�]� ���̡`�H$�QX�����U��`�H$�A\]�����������������U��`�P$�EP�EP�EPQ�J`�у�]� �����������̡`�H(�������U��`�H(�AV�u�R�Ѓ��    ^]��������������U��`�P(�R]����������������̡`�P(�B�����U��`�P(�R]�����������������U��`�P(�R]�����������������U��`�P(�R ]�����������������U��`�P(�E�RjP�EP��]� ��U��`�P(�E�R$P�EP�EP��]� �`�P(�B(����̡`�P(�B,����̡`�P(�B0�����U��`�P(�R4]�����������������U��`�P(�RX]�����������������U��`�P(�R\]�����������������U��`�P(�R`]�����������������U��`�P(�Rd]�����������������U��`�P(�Rh]�����������������U��`�P(�Rx]�����������������U��`�P(�Rl]�����������������U��`�P(�Rt]�����������������U��`�P(�Rp]�����������������U����`�E�    �E�    �P(�RhV�E�P���҅���   �E���uG�`�H�A�U�R�Ћ`�Q�E�RP�M�Q�ҡ`�H�A�U�R�Ѓ��   ^��]� �`�Qh�h8  P���   �Ћ`�����E��Q(u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P�fS����3�^��]� �M��U�j ���Q�MR�����E�P�<S�����   ^��]� �������������U��`��V��H�A�U�R�Ѓ��M�Q��������^u�`�B�P�M�Q�҃�3���]� �`�H$�E�I�U�RP�ы`�B�P�M�Q�҃��   ��]� �U��Q�`�P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U��`�P(�R8]�����������������U��`�P(�R<]�����������������U��`�P(�R@]�����������������U��`�P(�RD]�����������������U��`�P(�RH]�����������������U��`�P(�E�R|P�EP��]� ����U��`�P(�RL]�����������������U��`�E�P(�BT���$��]� ���U��`�E�P(�BPQ�$��]� ����̡`�H(�Q�����U��`�H(�AV�u�R�Ѓ��    ^]��������������U��`�P(���   ]��������������U��`�H(�A]����������������̡`�H,�Q,����̡`�P,�B4�����U��`�H,�A0V�u�R�Ѓ��    ^]�������������̡`�P,�B8�����U��`�P,�R<��VW�E�P�ҋu���`�H�QV�ҡ`�H$�QDV�ҡ`�H$�QLVW�ҡ`�H$�AH�U�R�Ћ`�Q�J�E�P�у�_��^��]� �������U��`�P,�E�R@��VWP�E�P�ҋu���`�H�QV�ҡ`�H�QVW�ҡ`�H�A�U�R�Ѓ�_��^��]� ��̡`�H,�j j �҃��������������U��`�P,�EP�EPQ�J�у�]� U��`�H,�AV�u�R�Ѓ��    ^]�������������̡`�P,�B����̡`�P,�B����̡`�P,�B����̡`�P,�B ����̡`�P,�B$����̡`�P,�B(�����U��`�P,�R]�����������������U��`�P,�R��VW�E�P�ҋu���`�H�QV�ҡ`�H$�QDV�ҡ`�H$�QLVW�ҡ`�H$�AH�U�R�Ћ`�Q�J�E�P�у�_��^��]� �������U��`�H��D  ]��������������U��`�H��H  ]��������������U��`�H��L  ]��������������U��`�H�I]�����������������U��`�H�A]�����������������U��`�H�I]�����������������U��`�H�A]�����������������U��`�H�I]�����������������U��`�H���  ]��������������U��`�H�A]�����������������U���V�u�E�P���k����`�Q$�J�E�P�у���u-�`�B$�PH�M�Q�ҡ`�H�A�U�R�Ѓ�3�^��]Ë`�Q�J�E�jP�у���u=�U�R��������u-�`�H$�AH�U�R�Ћ`�Q�J�E�P�у�3�^��]Ë`�B�HjV�у���u�`�B�HV�у����I����`�Q$�JH�E�P�ы`�B�P�M�Q�҃��   ^��]�����������U��`�H�A ]�����������������U��`�H�I(]�����������������U��`�H��  ]��������������U��`�H��   ]��������������U��`�H��  ]��������������U��`�H��  ]��������������U��`�H�A$��V�U�WR�Ћ`�Q�u���BV�Ћ`�Q$�BDV�Ћ`�Q$�BLVW�Ћ`�Q$�JH�E�P�ы`�B�P�M�Q�҃�_��^��]������U��`�H���  ��V�U�WR�Ћ`�Q�u���BV�Ћ`�Q$�BDV�Ћ`�Q$�BLVW�Ћ`�Q$�JH�E�P�ы`�B�P�M�Q�҃�_��^��]���U��`�H���  ]��������������U���<����SVW�E�    t�E�P�   �X������/�`�Q�J�E�P�   �ы`�B$�PD�M�Q�҃��}�`�H�u�QV�ҡ`�H$�QDV�ҡ`�H$�QLVW�҃���t)�`�H$�AH�U�R����Ћ`�Q�J�E�P�у���t&�`�B$�PH�M�Q�ҡ`�H�A�U�R�Ѓ�_��^[��]���U��`�H�U���  ��VWR�E�P�ы`�u���B�HV�ы`�B$�HDV�ы`�B$�HLVW�ы`�B$�PH�M�Q�ҡ`�H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]���������̡`�H���   ��U��`�H���   V�uV�҃��    ^]�������������U��`�P�]��`�P�B����̡`�P���   ��U��`�P�R`]�����������������U��`�P�Rd]�����������������U��`�P�Rh]�����������������U��`�P�Rl]�����������������U��`�P�Rp]�����������������U��`�P�Rt]�����������������U��`�P���   ]��������������U��`�P�Rx]�����������������U��`�P���   ]��������������U��`�P�R|]�����������������U��`�P���   ]��������������U��`�P���   ]��������������U��`�P���   ]��������������U��`�P���   ]��������������U��`�P���   ]��������������U��`�P���   ]��������������U��`�P���   ]��������������U��`�P���   ]��������������U��`�P���   ]��������������U��`�P���   ]��������������U��`�P�EPQ��  �у�]� �U��`�P���   ]��������������U��`�P���   ]��������������U��`�P���   ]��������������U��E��t �`�R P�B$Q�Ѓ���t	�   ]� 3�]� U��`�P �E�RLQ�MPQ�҃�]� U��E��u]� �`�R P�B(Q�Ѓ��   ]� ������U��`�P�R]�����������������U��`�P�R]�����������������U��`�P�R]�����������������U��`�P�R]�����������������U��`�P�R]�����������������U��`�P�R]�����������������U��`�P�E�R\P�EP��]� ����U��`�E�P�B ���$��]� ���U��`�E�P�B$Q�$��]� �����U��`�E�P�B(���$��]� ���U��`�P�R,]�����������������U��`�P�R0]�����������������U��`�P�R4]�����������������U��`�P�R8]�����������������U��`�P�R<]�����������������U��`�P�R@]�����������������U��`�P�RD]�����������������U��`�P�RH]�����������������U��`�P�RL]�����������������U��`�P�RP]�����������������U��`�P���   ]��������������U��`�P�RT]�����������������U��`�P�EPQ��  �у�]� �U��`�P���   ]��������������U��`�P���   ]��������������U��`�P�RX]����������������̡`�P���   ��U��`�P���   ]��������������U��`�P���   ]��������������U��`�P���   ]��������������U��`�P���   ]�������������̡`�P���   ��U��`�P���   ]�������������̡`�P���   ��`�P���   ��`�P���   ��U��`�H���   ]��������������U��`�H��   ]��������������U��`�H�U�E��VWRP���  �U�R�Ћ`�Q�u���BV�Ћ`�Q�BVW�Ћ`�Q�J�E�P�у�_��^��]������������U��`�H���  ]��������������U��`�} �P(�R8��P��]� ����U��`�P�BdS�]VW��j ���Ћ`�Q�����   h���hc  V�Ћ`�����Eu�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћ`�Q(�BHV���Ѕ�t �`�Q(�E�R VP���҅�t�   �3��EP�p>����_��^[]� ����U���V�E���MP�{���P���#����`�Q�J���E�P�у���^��]� ��̡`�PD�BQ�Ѓ���������������̡`�PD�BQ�Ѓ���������������̡`�PD�BQ�Ѓ����������������U��`�PX��Q�
�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ���������U��`�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U��`�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U��`�PX��`VWQ�J�E�P�ы��E���   ���_^��]� �������������U��`�PX�EPQ�J�у�]� ����U��`�PX�EPQ�J�у�]� ����U��`�PX�EPQ�J�у�]� ����U��`�PX�EPQ�J�у�]� ����U��`�PX�EPQ�J$�у�]� ����U��`�PX�EPQ�J �у�]� ����U��`�PD�EP�EPQ�J�у�]� U��`�HD�U�j R�Ѓ�]�������U��`�H@�AV�u�R�Ѓ��    ^]��������������U��`�HD�	]��U��`�H@�AV�u�R�Ѓ��    ^]��������������U��`�HD�U�j R�Ѓ�]�������U��`�H@�AV�u�R�Ѓ��    ^]��������������U��`�U�HD�Rh'  �Ѓ�]����U��`�H@�AV�u�R�Ѓ��    ^]�������������̡`�HD�j h�  �҃�����������U��`�H@�AV�u�R�Ѓ��    ^]�������������̡`�HD�j h:  �҃�����������U��`�H@�AV�u�R�Ѓ��    ^]��������������U���3��E��E��`���   �R�E�Pj�����#E���]�̡`�HD�j h�F �҃�����������U��`�H@�AV�u�R�Ѓ��    ^]�������������̡`�HD�j h�_ �҃�����������U��`�H@�AV�u�R�Ѓ��    ^]��������������U��E����u��]� �E��`�E�    ���   �R�E�Pj������؋�]� ̡`�PD�B$Q�Ѓ���������������̡`�PD�B(Q�Ѓ���������������̡`�PD�BQ�Ѓ���������������̡`�PD�B(Q�Ѓ���������������̡`�PD�BQ�Ѓ���������������̡`�PD�B(Q�Ѓ���������������̡`�PD�BQ�Ѓ���������������̡`�PD�B(Q�Ѓ���������������̡`�PD�BQ�Ѓ���������������̡`�PD�B(Q�Ѓ���������������̡`�PD�BQ�Ѓ���������������̡`�PD�B(Q�Ѓ���������������̡`�PD�BQ�Ѓ���������������̡`�PD�B(Q�Ѓ���������������̡`�PD�BQ�Ѓ���������������̡`�PD�B(Q�Ѓ���������������̡`�PD�BQ�Ѓ���������������̡`�PD�B(Q�Ѓ���������������̡`�PD�BQ�Ѓ����������������U��M�EV�u������t#W���    �Pf�y������f�8f�u�_^]� �U��� �E���M��"  �ȉES���V�u��W�}�ǃ��Q���ƃ��։E��B��E���؉M�E��U���M��~�U�U���)}�M��>���E��}�t�u+���I �\�P���m���u�E�����E��   )}��u��	;]��u��s���u;]�]�}�M��>P�E�V�Ѕ�}	�u���]�M��E��VP�҅��V������F��}�t!�M�+ȃ����\�P���m���u�]��;]~�����_^[��]� ���U���(W�}�����E�E���M��  �MS�؉E������ǃ��S�����E�ы���V�]�U��E܉U���]��~�E�E��)}��]��)�M�U��E�Q�M�RP������E�����E��   )}��u�;E��؉u�s���u;]�]�}�M���>P�E؋V�Ѕ�}	�u؃��]��M���E�VP�҅��i����}���F�t&�M�+ȃ���I �Pf�\����f�f�u�]��}�;E�w����%���^[_��]� ��������U���(W�}�����E�E���M��)  �ЉE������ǃ��J���SV�uƃ��ΉE��A��E����؉U��E܉M����I �U���~�M�M��)}��U��A�M�ɋE��M�t�M�+���I �\�p���m���4u�E�����E��   )}��u�;E��؉u�s���u;]�]�}�M��>P�E؋V�Ѕ�}	�u؃��]��M��E�VP�҅��Q����}���F�t�M�+ȃ���\�P������u�]��}�;E~�����^[_��]� ���������������U��E�Pu�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����E��SV��W�]�t8�u��t1�}��t*�} t$�VP��Ѕ���   |������E�   �}}_^3�[��]� �}�M���E�������uu��VP�҅�t#}����}����}��E9E�~�_^3�[��]� ��~3�E���]��]�E��E�M���؋ESP���҅�u�����_��^[��]� ���������������U����E��SV��W�]��  �u����   �}����   �} ��   �VP��Ѕ���   }�M_^�    3�[��]� �O�3����E�   �M} ����   �E���8_^3�[��]� ���M�U���<�M������uuVQ���҅�t}�O��M��W�U��M9M�~�뤅�~3�E���]��]�E��E�M���؋ESP���҅�u�����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� �����������U��V�u�F��F�����������������ܛ  ����������D�Ez��^�P�P�]��������������N�X�N^�X]�������P�P��P(�P �P�P@�P8�P0�PX�PP�PH����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX��������U��M�A8��   �IXV�AP�I@���I�AP�I(�AX�I ���I0���A@�I �A8�I(���IH����������Dz�u�؋��5�����^��]���W���A�IX�AP�I�A8�I�A�I@�AP�I@�U��A8�IX�]������IH�����I0�����e��	����ݝx����A�I(�U��A�I �U��AX�I �]��AP�I(�����IH�E����	���������I�������]��A8�I(�A@�I �����	�������I���E��e��I0�������]��E��e����]����e��ˋE��x������]������]��AH�I@�A0�IX�����]��AX�I�AH�I(�����]��A0�I(�A@�I�����]��AP�I0�AH�I8�����]��AH�I �AP�I�����]��A8�I�A0�I �   �����]��_^��]�������U��y0 ts��U�����Au���A�Z����Au�B�Y�A�Z����Au�B�Y�A�����z��Y�A �Z����z�B�Y �A(�Z����zZ�B�Y(]� �E��Q�P�Q�P�Q �P�Q$�P�Q(�@�A,�Q�A��Q �A�A$�Q�Q(�A�A,�Q�A�A0   ]� U��y0 tL��E�A�A �A�A(�A�0�����������X�X�A� �A �`�A(�`�E����X�X]� ��E����������P���P�E����X�X]� ��̋�3ɉ�H�H�H�V��V��+���FP�+��3����F�F^��3���A�A�A����A�`�
�@�b�	���B�a�������U����   ��UV���q�U�W3��<��M��}���  ��S�]�k  ��؋�U��M�U��U�@�����@�U��@�B�@�������@���@�G�>��w����U���  �w������݃��B��   �U������ɋP��R�э����]��B���B�P���R���U����E������]��E��M��E������������]��E����E����E��E��]����E��]����E��]��]����U��E��U�����B���B���U������������]��E����E����������E������E��E��]����E��]����E��]����U��E��]���R�э�������B���B�P���R���U����E��������]��E����E����������E������E��E��]��E��]����E��]��U��E��]�����B���B���U����E��������]��E����E����������E������E��E��]��E��]����E��]��E��U��`�����E�U���������;���   �ލ�+���͋�@����������]��@���]��@���U������M������]��E��E����E��������]��E������������E��E��]��E��E��]����E��]��E��U�u�������������������������������M���Q�ʍU��R���[�[������E�KH��P�E��SL��H�щKP�P�ST�H�KX�P�������S\z^�E�����������zP���CP�����CX���CH���CX�������cH���[�[ �[(�C(�KP�C �KX���C�KX�C(�KH���CH�K �\���E���������za�CX�����CP�����cH�CH���CP�������[���[ �[(�CP�K(�C �KX���C�KX�CH�K(���C �KH�C�KP�����[0�[8�[@�[�CP�����CX�����KH�CX�����cP���[0�[8�[@�C8�KX�C@�KP���C@�KH�CX�K0���CP�K0�C8�KH�����[�[ �[(��$���SP������E��U�   �����}��M�����م�~�A8����u��1���U�@���K�I��@�K0���CH�H��� �K �C�@�K8���@�KP���C(��C�@�K@���CX�H�D��@�����U���]��C���@�K0���CH�H���C ��C�@�K8���@�KP���C(��C�C@�H���CX�H3������U��x  �A������܃��E����E   �E�
���������ɋE������׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H�E������������������������������E����]��E��]����]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H�E��������]������M������������������������]��E��]��E��]�׋��@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H���]������M������������������������]��E�Eȃ��]���E����]ȃE׃m����@�E�Ѝ��K��@�K0���CH�H��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H���]������M������������������������U��E��]��E��U�������E������������;���   �P�U��+ЉU�
���������ʋE���׋��U�@���K��@�K0���CH�H���]�� �K �C�@�K8���@�KP���]�� �K(�C�C@�H���CX�H�   E)E���]����E��������������������M����������]��E��E��U�����[������_��^��]� ��[��_��^���؋�]� �����������hxPh_� ��G  ���������������hxjh_� �G  ����uË@����U��V�u�> t/hxjh_� �G  ����t��U�M�@R�Ѓ��    ^]���U��Vhxjh_� ���IG  ����t�@��t�MQ����^]� 3�^]� �������U��Vhxjh_� ���	G  ����t�@��t�MQ����^]� 3�^]� �������U��Vhxjh_� ����F  ����t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vhxjh_� ���yF  ����t�@��t�MQ����^]� 3�^]� �������U��Vhxj h_� ���9F  ����t�@ ��t�MQ����^]� 3�^]� �������U��Vhxj$h_� ����E  ����t�@$��t�MQ����^]� 2�^]� �������Vhxj(h_� ���E  ����t�@(��t��^��3�^������Vhxj,h_� ���E  ����t�@,��t��^��3�^������U��Vhxj0h_� ���YE  ����t�@0��t�MQ����^]� 3�^]� �������U��Vhxj4h_� ���E  ����t�@4��t�M�UQR����^]� ���^]� ��Vhxj8h_� ����D  ����t�@8��t��^��3�^������U��Vhxj<h_� ���D  ����t�@<��t�MQ����^]� ��������������U��Vhxj@h_� ���iD  ����t�@@��t�MQ����^]� ��������������U��VhxjDh_� ���)D  ����t�@D��t�MQ����^]� 3�^]� �������U��VhxjHh_� ����C  ����t�@H��t�MQ����^]� ��������������VhxjLh_� ���C  ����t�@L��t��^��3�^������VhxjPh_� ���|C  ����t�@P��t��^��3�^������VhxjTh_� ���LC  ����t�@T��t��^��^��������VhxjXh_� ���C  ����t�@X��t��^��^��������Vhxj\h_� ����B  ����t�@\��t��^��^��������U��Vhxj`h_� ���B  ����t�@`��t�M�UQR����^]� 3�^]� ���U��Vhxjdh_� ���yB  ����t�@d��t�M�UQR����^]� 3�^]� ���U��Vhxjhh_� ���9B  ����t�@h��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vhxjlh_� ����A  ����t�@l��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vhxjph_� ���A  ����t�@p��t�M�UQR����^]� 3�^]� ���U��Vhxjth_� ���YA  ����t�@t��t�M�UQR����^]� 3�^]� ���U��Vhxjxh_� ���A  ����t�@x��t�M�UQR����^]� 3�^]� ���U��Vhxj|h_� ����@  ����t�@|��t�MQ����^]� 3�^]� �������U��Vhxh�   h_� ���@  ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vhxh�   h_� ���F@  ����t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vhxh�   h_� ����?  ����t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vhxh�   h_� ���?  ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U���|��A�����U����U����U��  S�V�E��EW�����������   ���������U�r�z�
�R;��4v���4��I�$ȍ��F�R�a���F�a�uB�!�]��B�a�U��B�a�U������������]��E����E����������E��������E��G��$ȍ��]��B�a�U��B�a�U������������]��E����E����������E��������E��������m�������_�U�^��[�U����U����������������������  ����������D�Ez���P�P���]� �������E�����E����X�M��X��]� �������U���@�(��A�������E�    ���]����]��]�� ��������]����]��]���   �	S�]VW�M��E����������t[��%�����E�M�����@��P������F�@��R�M������~���Q�M������v;�t�v��P�M������M����m��M�u�_^[�M�UQR�M��A�����]� ����������̋Q3���|�	��t��~�    t������u��3�������U��QV�u;��}�	���    u����;�|���^]� +ƃ�^]� �������U��VW�}��|-�1��t'�Q3���~�΍I �1�������;�t����;�|���_^]� �������������̋Q3���~%V�1�d$ ���   @u�����t������u�^�̋QV3���~�	�d$ ����Шt������u��^�������U��Q3�9A~��I ��$��������;A|�Q��~[SVW�   3ۋ���x5��%���;��E���}$��������%���;E�u�
   ���;q|݋Q���G���;�|�_^[��]�������U��	����%�����E��   @t����������wg�$��Z�E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� 4ZJZ]ZqZ�Z����U����S��V������   @Wt���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V��V����FP���3����F�F^��U��SV��WV�r���^S�i���E3���;ǉ~�~t_�`�Q���   h8���jIP�у�;ǉt9�}��t;�`�B���   h8���    jNQ�҃����uV������_^3�[]� �E�~_�F^�   []� ����������U��SV��WV�����^S����}3Ƀ�;��N�N��   9��   �G;���   �`�Q���  h8���jlP�у����t=� t@�G��t9�`�Jh8���    ���  jqR�Ѓ����u���]���_^3�[]� �O�N�G�Q��    R�F�QP�  �����t�N�WP��QPR�h  ��_^�   []� ���������U��SV��WV�����~W���3Ƀ�9M�N�N��   �E;���   ��    �`�H���  h8�h�   S�҃����t=�} tH�E��tA�`�Q���  h8���h�   P�у����u���b���_^3�[]� �U�V�,�F   �`�H���  h8�h�   j�҃����t��E�M�F�PSPQ�a  �E����t!�V�?�W�RWP�E  ��_^�   []� ��M�_^�   []� ���U��Q2���~CS�]V�1W������������;�u��   @u�����u3���   ��
���u�_^[��]� �����������U��S�]V��3�W�~���F�F�C;CV��   ���W���3��F�F�`�Q���   h8�jIj�Ѓ������   �`�Q���   h8�jNj�Ѓ����uV�����_��^[]� ��F   �F   ����K�H�C��B�_��^�   []� �p��W�j��3��F�F�`�B���   h8�jIj�у����t[�`�B���   h8�jNj�у�����\�����F   �F   ����S�Q��K�H��C�B��   _��^[]� �����������U��3�V���F�F�F�EP�������^]� �������������U��EVP���������^]� ����������U��U��t�M��t�E��tPRQ�s  ��]�����������̡`�H���   ��U��`�H���   V�u�R�Ѓ��    ^]����������̡`�P���   Q�Ѓ�������������U��`�P�EPQ���   �у�]� ̡`�H�������U��`�H�AV�u�R�Ѓ��    ^]��������������U��`�H�AV�u�R�Ѓ��    ^]��������������U��`�P��Vh�  Q���   �E�P�ы`���   �Q8P�ҋ�`���   ��U�R�Ѓ���^��]��������������̡`�P�BQ�Ѓ����������������U��`�P�EPQ�J\�у�]� ����U��`�P�EP�EP�EP�EP�EPQ���   �у�]� �U��`�P�EP�EP�EP�EPQ�JX�у�]� �������̡`�P�B Q��Y�U��`�P�EP�EP�EP�EPQ���   �у�]� �����U��`�P�EP�EP�EPQ�J�у�]� ������������U��`�H��   ]��������������U��`�P�R$]�����������������U��`�P�EP�EP�EP�EPQ�J(�у�]� ��������U��`�P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U��`�P�EP�EP�EP�EPQ�J,�у�]� ��������U��`V��H�QWV�ҋ��`�H�QV�ҋ`�Q�M�R4Q�MQ�MQ���W���Pj j V�҃�(_^]� �����������U��`�P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U��`�P�EP�EPQ�J@�у�]� U��`�P�EPQ�JD�у�]� ���̡`�P�BLQ�Ѓ���������������̡`�P�BLQ�Ѓ���������������̡`�P�BPQ�Ѓ����������������U��`�P�EPQ�JT�у�]� ����U��`�P�EPQ�JT�у�]� ����U��`�P�EP�EPQ���   �у�]� �������������U��`�P�E���   ��VP�EPQ�M�Q�ҋu�    �F    �`���   j P�BV�Ћ`���   �
�E�P�у� ��^��]� ������̡`�P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡`�H�������U��`�H�AV�u�R�Ѓ��    ^]��������������U��`�P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U��`�P�EPQ�J�у�]� ���̡`�P�BQ��Y�U��`�P�EP�EPQ�J�у�]� U��VW�������M�U�x@�EPQR������H ���_^]� �U��VW������M�U�xD�EPQR������H ���_^]� �V���x���xH u3�^�W���f���΍xH�\���H �_^�����U��V���E���xL u3�^]� W���0���M�U�xL�EPQR������H ���_^]� �������������U��V�������xP u���^]� W�������M�U�xP�EP�EQRP�������H ���_^]� ��������U��V������xT u���^]� W������M�xT�EPQ���}���H ���_^]� U���S�]��VW��t.�M�薃�����O���xL�E�P���A���H ��ҍM��Ѓ���}��tZ�`�H�A�U�R�Ћ`�Q�J�E�WP�ы`�B�P�M�Q�҃��������@@��t�`�QWP�B�Ѓ�_^[��]� ������U��VW������xH�EP������H ���_^]� ���������U��VW������M�U�xD�EP�EQRP���j���H ���_^]� �������������U��V���E���xP u
�����^]� W���-���M�U�xP�EP�EQ�MR�UPQR������H ���_^]� ��������������U��V���� ���xT u
�����^]� W���� ���M�xT�EPQ��� ���H ���_^]� ��������������U��V��� ���xX tW��� ���xX�EP���y ���H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u��O  ����t.�E�;�t'�`�J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡`�H��   ��U��`�H��$  V�u�R�Ѓ��    ^]�����������U��`�UV��H��(  VR�Ѓ���^]� �����������U��`�P�EQ��,  P�у�]� �U��`�P�EQ��,  P�у������]� ���������̡`�H��0  ��`�H��4  ��U��E��t�@�3��`�RP��8  Q�Ѓ�]� �����U��`�P�EPQ��<  �у�]� �U��`�P�EP�EP�EPQ��@  �у�]� ���������U��`�P�EP�EPQ��D  �у�]� �������������U��`�P�EPQ��H  �у�]� �U��`�P�E��L  ��VWPQ�M�Q�ҋu���`�H�QV�ҡ`�H�QVW�ҡ`�H�A�U�R�Ѓ�_��^��]� ��������������̡`�P��T  Q�Ѓ������������̡`�P��P  Q�Ѓ�������������U��`�P�EPQ��X  �у�]� ̡`�H��\  ��U��`�H��`  V�u�R�Ѓ��    ^]�����������U��`�P�EP�EP�EP�EP�EPQ��d  �у�]� �U��`�P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���w��������3��F�F �F$�F(�F,�F0�F4�F8�F<�F@�FD�FH�FL�FP�FT�FX�_p��G`�Gd�Gh�Gx�����G|   ��_^��������������V��W�>��t7���O����xP t$S���A���j j �XPj�FP���-����H ���[�    �~` t�`�H�V`�AR�Ѓ��F`    _^������������U��SV��Fx�`�Q��   WV�^dSP�EP�~`W�у����F|��   �> ��   �; ��   �U�~pW�^hSR�ļ������u#���h���`�H��0  h�   �҃��E�~P��輧���j j jW�N������F|t��������F|_^[]� �F|_�Fx����^[]� �F|�����    �`�Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��V��~d �F`tLW�};~xtBWPj�NQ��������F|u�E���~xt�    �F`_^]� �M���Fx����t�3�_^]� U��QVW�}����L  �`�H�QhV�҃����`u"�H��0  h��h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���t�3�9u�~!�E���<� t��Q����I  �E��;u�|�UR�{�����_�   ^��]� �����������U��QVW�}����NK  �`�H�QhV�҃����`u"�H��0  h��h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���tЋE��t�3�9u�~:��E�<� t'���`�QP�Bh�Ѓ���t�M��R����H  ��;u�|ȍEP������_�   ^��]� �����������h��h�   h�h�   �g������t�������3��������V���(����N^鯡�����������������U��VW�}�7��t��������N胡��V�M �����    _^]�U���EV���V��������Au�`�H��0  hжj,�����^��^]� �����U���W������G���U����������A�  ������A��   � �������AuR������AuKV����_  ����_  �ȅ�u��^����__��]Ëƙ����ҋ�u�u��E�^������__��]���������Au������=���������Au6�����������U������G�����_��������Au�����U����_�
����������h  �E����U��0���������A{���������__��]�������������__��]����U���0�V�E��������At���(�������Au������H����0��$�
e  ����H����^�e�����^]� ��������������U����V�E��������u�   �3����]����Az�   �3�3����0�;���W���$���d  ��E���0��$�|d  �V����������Au�`�H��0  hжj�����^����_u������������^]� ���U������EV�ы�������z!�`�؋H��0  hжj5�����U������$��c  �]��F�$��c  �}��$��c  ��E�$��c  �^�����&���^��]� ���������������U��`���   �BXQ�Ѓ���u]� �`�Q|�M�RQ�MQP�҃�]� ���U��`���   �BXQ�Ѓ���u]� �`�Q|�M�R8Q�MQP�҃�]� ���U��EV��j ��`�Qj j P�B�ЉF����^]� ��̡`Vj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� �`�Q�MP�EP�Q�JP�у��F�   ^]� ����U��M��P]����U��M��P]����U��M��P]����V���<��F    �`�HP�hPwVh@wh0w�҉F����^����������̃y �<�u�`�PP�A�JP��Y��U��A��u]� �`�QP�M�Rj Q�MQP�҃�]� ��U��A��t�`�QP�M�RQP�҃�]� ������������U��A��t�`�QP�M�RQP�҃�]� �����������̡`�HP���   ��U��`�HP���   ]�������������̡`�HP�QP�����U��`�HP�AT]����������������̋��     �@    �V����t)�`�QPP�BL�Ћ`�QP��J<P�у��    ^�������������U��SV�ً3�;�Wt�`�QPP�B<�Ѓ��3�s�}�EhPwW�C�`�QP�J8h@wh0wP�EP�у�9u�~O�I ���z u!���@   �`�QP���H�RQ�҃��`�HP��A@VR�Ћ�����;u�A|�3�9_^��[]� ������U��SVW��3�9w~>�]�`�HP��A@VR�Ѓ���t/�`�QPj SjP�B�Ѓ���t��;w|�_^�   []� �`�QP��JLP�у�_^3�[]� ���������̡`�PP��JDP�у�������������̡`�PP��JHP��Y��������������̡`�PP��JLP��Y���������������U��U�E�@R�URP�I���]� �����3���������������U��V��~ �<�u�`�HP�V�AR�Ѓ��Et	V��������^]� ����h|PhD �   ���������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d��������]� ���������U��h|jhD �,  ����t
�@��t]��3�]��������Vh|j\hD ����  ����t�@\��tV�Ѓ���^�����Vh|j`hD ����  ����t�@`��tV�Ѓ�^�������U��Vh|jdhD ���  ����t�@d��t
�MQV�Ѓ�^]� ������������U��Vh|jhhD ���Y  ����t�@h��t
�MQV�Ѓ�^]� ������������Vh|jlhD ���  ����t�@l��tV�Ѓ�^�������U��Vh|h�   hD ����  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh|h�   hD ���  ����t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh|jphD ���I  ����t�@p��t�MQV�Ѓ�^]� ��^]� ��U��Vh|jxhD ���	  ����t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh|jxhD ����  ����t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh|jxhD ���  ����t�@|��t�MVQ�Ѓ������^]� �   ^]� ����������̋���������������h|jhD �/  ����t	�@��t��3��������������U��V�u�> t+h|jhD ��  ����t�@��tV�Ѓ��    ^]�������U��VW�}����t0h|jhD �  ����t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh|jhD ���i  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh|jhD ���)  ����t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh|j hD ����  ����t�@ ��tV�Ѓ�^�3�^���Vh|j$hD ���  ����t�@$��tV�Ѓ�^�3�^���U��Vh|j(hD ���  ����t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh|j,hD ���9  ����t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh|j(hD ����  ����t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh|j4hD ���  ����t�@4��tV�Ѓ�^�3�^���U��Vh|j8hD ���y  ����t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh|j<hD ���)  ����t�@<��t
�MQV�Ѓ�^]� ������������Vh|jDhD ����  ����t�@D��tV�Ѓ�^�3�^���U��Vh|jHhD ���  ����t�M�PHQV�҃�^]� U��Vh|jLhD ���  ����u^]� �M�PLQV�҃�^]� �����������U��Vh|jPhD ���I  ����u^]� �M�U�@PQRV�Ѓ�^]� �������Vh|jThD ���  ����u^Ë@TV�Ѓ�^���������U��Vh|jXhD ����  ����t�M�PXQV�҃�^]� U��Vh|h�   hD ���  ����u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh|h�   hD ���V  ����u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh|h�   hD ���  ����u^]� �M���   QV�҃�^]� �����U��Vh|h�   hD ����  ����u^]� �M���   QV�҃�^]� �����U��Vh|h�   hD ���  ����u^]� �M���   QV�҃�^]� �����U��Vh|h�   hD ���F  ����t�M�UQ�MR���   QV�҃�^]� ��U���Vh|h�   hD �  ����u�`�H�u�QV�҃���^��]ËM���   WQ�U�R�Ћ`�Q�u���BV�Ћ`�Q�BVW�Ћ`�Q�J�E�P�у�_��^��]��U��Vh|h�   hD ���v  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh|h�   hD ���&  ����t���   ��t�MQ����^]� 3�^]� �U��Vh|h�   hD ����  ����t���   ��t�MQ����^]� 3�^]� �U��Vh|h�   hD ���  ����t���   ��t�MQ����^]� 3�^]� �Vh|h�   hD ���i  ����t���   ��t��^��3�^����������������U��Vh|h�   hD ���&  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh|h�   hD ����  ����t���   ��t�MQ����^]� ��������U��Vh|h�   hD ���  ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vh|h�   hD ���I  ����t���   ��t��^��3�^����������������VW��3����$    �h|jphD ��  ����t�@p��t	VW�Ѓ�����8 t����_��^�����U��SW��3�V��    h|jphD �  ����t�@p��t	WS�Ѓ�����8 tsh|jphD �}  ����t�@p��t�MWQ�Ѓ������h|jphD �K  ����t�@p��t	WS�Ѓ����V���7�����t���[����E��^t�8��~=h|jphD ��  ����t�@p��t	WS�Ѓ�����8 u_�   []� _3�[]� ��������U��Vh|j\hD ���  ����t3�@\��t,V��h|jxhD �  ����t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh|j\hD ���I  ����t3�@\��t,V��h|jdhD �'  ����t�@d��t
�MQV�Ѓ���^]� ��������U���Vh|j\hD ����
  ����tG�@\��t@V�ЋEh|jdhD �E��E�    �E�    �
  ����t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh|j\hD ���i
  ����t\�@\��tUV��h|jdhD �G
  ����t�@d��t
�MQV�Ѓ�h|jhhD �
  ����t�@h��t
�URV�Ѓ���^]� ���������������U��Vh|j\hD ����	  ������   �@\��t~V��h|jdhD �	  ����t�@d��t
�MQV�Ѓ�h|jhhD �	  ����t�@h��t
�URV�Ѓ�h|jhhD �a	  ����t�@h��t
�MQV�Ѓ���^]� ��U���Vh|jthD ���&	  ����tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h|j`hD ��  ����t(�@`��t!�M�Q�Ѓ���^��]� �uh����_�����^��]� ������U���Vh|h�   hD ���  ����tR���   ��tH�MQ�U�R���ЋuP������h|j`hD �Z  ����t<�@`��t5�M�Q�Ѓ���^��]� �u�U�R���E�    �E�    �E�    ������^��]� �������������̋�3ɉH��H�@   �������������U��ыM��tK�E��t�`���   P�B@��]� �E��t�`���   P�BD��]� �`���   R�PD��]� �����U��`�P@�Rd]�����������������U��`�P@�Rh]�����������������U��`�P@�Rl]�����������������U��`�P@�Rp]�����������������U��`���   ���   ]�����������U��`���   ���   ]����������̡`�P@�Bt����̡`�P@�Bx�����U��`�P@�R|]����������������̡`�P@���   ��`���   �Bt��U��`�P@���   ]�������������̡`�P@���   ��U��`�P@���   ]��������������U��`�P@���   ]��������������U��`�P@���   ]��������������U��`�P@���   ]��������������U��`V��H@�QV�ҋM����t��#����`�Q@P�BV�Ѓ�^]� �̡`�PH���   Q�Ѓ�������������U��`�P@�EPQ�JL�у�]� ���̡`�P@�BHQ�Ѓ����������������U��`�P@�EP�EP�EPQ�J�у�]� ������������U��`�P@�EPQ�J�у�]� ����U��`�P@�EP�EPQ�J�у�]� U��`�P@�EPQ�J �у�]� ����U��`���   �R]��������������U��`���   �R]��������������U��`���   �R ]��������������U��`���   ���   ]�����������U��`���   ��D  ]�����������U��`�E���   �E ���   P�E���$P�EP�EP�EP��]� ���������U��`���   ���   ]����������̡`���   �B$��`�H@�Q0�����U��`�H@�A4j�URj �Ѓ�]����U��`�H@�A4j�URh   @�Ѓ�]�U��`�H@�U�E�I4RPj �у�]�̡`�H|�������U��V�u���t�`�Q|P�B�Ѓ��    ^]��������̡`�H|�Q �����U��V�u���t�`�Q|P�B(�Ѓ��    ^]��������̡`�H@�Q0�����U��V�u���t�`�Q@P�B�Ѓ��    ^]���������U��`�H@���   ]��������������U��V�u���t�`�Q@P�B�Ѓ��    ^]��������̡`�PH���   Q�Ѓ�������������U��`�PH�EPQ��d  �у�]� �U��`�H �IH]�����������������U��}qF uHV�u��t?�`���   �BDW�}W���Ћ`�Q@�B,W�Ћ`�Q�M�Rp��VQ����_^]����������̡`�P@�BT�����U��`�P@�RX]�����������������U��`�P@�R\]����������������̡`�P@�B`�����U��`�H��T  ]��������������U��`�H@�U�A,SVWR�Ћ`�Q@�J,���EP�ы`�Z��h��hE  �΋��&Y��Ph��hE  ���Y��P��T  �Ѓ�_^[]����U��E�M�UP��P�EjP�s�����]��������������̸   �����������U��V�u��t���u8�EjP�t�������u3�^]Ë��a�����t���t��U3�;P����#�^]�����h�Ph^� �������������������U��Vh�jh^� ���y�������t�@��t�M�UQRV�Ѓ�^]� 3�^]� �Vh�jh^� ���<�������t�@��tV�Ѓ�^�3�^���U��Vh�jh^� ���	�������t�@��t�M�UQRV�Ѓ�^]� ���^]� U���  Vh�jh^� �����������t/�@��t(�MWQ��x���VR�Ћ��E���b   ���_^��]� �u���ө���N`�˩�����   �������   赩����ݞ�  ��^��]� ����U��Vh�jh^� ���9�������t�@��t�M�UQRV�Ѓ�^]� ��������U��Vh�jh^� �����������t�@��t�M�UQ�MRQV�Ѓ�^]� ����U��Vh�j h^� ����������t�@ ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh�j$h^� ���i�������t�@$��t�MQV�Ѓ�^]� 3�^]� �����U��Vh�j(h^� ���)�������t�@(��t�M�UQ�MR�UQRV�Ѓ�^]� U��QVh�j,h^� �����������t �@,���E�t�E�MPQV�U���^��]� ��^��]� ��������U��Vh�j0h^� ����������t#�@0��t�E�M�U���$QRV�Ѓ�^]� 3�^]� ��������Vh�j4h^� ���L�������t�@4��tV�Ѓ�^�3�^���Vh�j8h^� ����������t�@8��tV�Ѓ�^�������U���`Vh�jDh^� �����������t(�@D��t!W�M�VQ�Ћ��E���   ���_^��]� �u���������^��]� ����U��Vh�jHh^� ����������t�@H��t
�MQV�Ѓ�^]� ������������U��Vh�jLh^� ���I�������t�@L��t�MQV�Ѓ�^]� ���^]� ����U��Vh�jPh^� ���	�������t�@P��t
�MQV�Ѓ�^]� ������������U��Vh�jTh^� �����������t�@T��t
�MQV�Ѓ�^]� ������������U��Vh�jXh^� ����������t.�@X��t'�M �UQ�MR�UQ�MR�UQ�MRQV�Ѓ� ^]� 3�^]� �������������Vh�j`h^� ���,�������t�@`��tV�Ѓ�^�3�^���U��Vh�jdh^� �����������t�@d��t�MQV�Ѓ�^]� 3�^]� �����U���Vh�jhh^� ����������t1�@h��t*�MQ�U�VR�Ћu��P��������M�������^��]� �u���d�����^��]� �����������Vh�jph^� ���L�������t�@p��tV�Ѓ�^Ã��^��Vh�jlh^� ����������t�@l��tV�Ѓ�^Ã��^��Vh�jth^� �����������t�@t��tV�Ѓ�^�3�^���U��Vh�jxh^� ����������t�@x��t
�MQV�Ѓ�^]� ������������Vh�j|h^� ���|�������t�@|��tV�Ѓ�^�������Vh�h�   h^� ���I�������t���   ��tV�Ѓ�^�U��Vh�h�   h^� ����������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������U��Vh�h�   h^� �����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U���Vh�h�   h^� ���s�������tU���   ��tKW�M�VQ�Ћ`�u���B�HV�ы`�B�HVW�ы`�B�P�M�Q�҃�_��^��]� �`�H�u�QV�҃���^��]� ����������Vh�h�   h^� �����������t���   ��tV�Ѓ�^Ã��^������������U��Vh�h�   h^� ����������t���   ��t
�MQV�Ѓ�^]� ������U��Vh�h�   h^� ���V�������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������Vh�h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������U��Vh�h�   h^� ���v�������t%���   ��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���U��Vh�h�   h^� ���&�������t���   ��t�M�UQRV�Ѓ�^]� ���^]� ����������U��Vh�h�   h^� �����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�h�   h^� ����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�h�   h^� ���6�������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�h�   h^� �����������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������Vh�h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������Vh�h�   h^� ���Y�������t���   ��tV�Ѓ�^�3�^�������������Vh�h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������Vh�h�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������U��Vh�h�   h^� ����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������Vh�h�   h^� ���I�������t���   ��tV�Ѓ�^�3�^�������������U���Vh�h�   h^� ����������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh�h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ��Vh�h�   h^� ���I�������t���   ��tV�Ѓ�^�3�^�������������U���Vh�h�   h^� ����������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh�h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ��Vh�h�   h^� ���I�������t���   ��tV�Ѓ�^�3�^�������������U��Vh�h�   h^� ����������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��QVh�h�   h^� ����������t#���   ���E�t�E�MPQV�U���^��]� ��^��]� ��U��Vh�h�   h^� ���f�������t!���   ��t�E�M�U���$QRV�Ѓ�^]� ���������U��Vh�h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�h�   h^� �����������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�h   h^� ���v�������t��   ��t�MQV�Ѓ�^]� 3�^]� ���������������Vh�h  h^� ���)�������t��  ��tV�Ѓ�^�3�^�������������U���Vh�h  h^� �����������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh�h  h^� ���c�������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh�h  h^� �����������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U��Vh�h  h^� ���f�������t��  ��t
�MQV�Ѓ�^]� ������U��Vh�h  h^� ���&�������t��  ��t
�MQV�Ѓ�^]� ������U��Vh�h  h^� �����������t��  ��t
�MQV�Ѓ�^]� ������Vh�h   h^� ����������t��   ��tV�Ѓ�^�3�^�������������U��Vh�h$  h^� ���f�������t��$  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�h(  h^� ����������t!��(  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�h,  h^� �����������t��,  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh�h0  h^� ���y�������t��0  ��tV�Ѓ�^�3�^�������������U��Vh�h4  h^� ���6�������t��4  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�h8  h^� �����������t��8  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�h<  h^� ����������t��<  ��t�M�UQ�MRQV�Ѓ�^]� ��������������U��Vh�h@  h^� ���F�������t��@  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh�hD  h^� �����������t��D  ��tV�Ѓ�^�3�^�������������U��Vh�hH  h^� ����������t��H  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�hL  h^� ���f�������t��L  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�hP  h^� ����������t!��P  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��QVh�hT  h^� �����������t'��T  ���E�t�E�M�UPQRV�U���^��]� ��^��]� ��������������U��Vh�hX  h^� ���f�������t%��X  ��t�E�M�U���$Q�MRQV�Ѓ�^]� �����U��Vh�j<h^� ����������t�@<��t�M�UQRV�Ѓ�^]� ��������U��Vh�j@h^� �����������t�@@��t�MQV�Ѓ�^]� 3�^]� �����h�Ph�� �������������������h�jh�� ��������uË@����U��V�u�> t/h�jh�� �S�������t��U�M�@R�Ѓ��    ^]���U��Vh�jh�� ����������t �@��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�jh�� �����������t�@��t�M�UQR����^]� ����������U��Vh�jh�� ����������t�@��t�M�UQR����^]� ����������U��Vh�jh�� ���I�������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh�j h�� �����������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh�j$h�� ����������t �@$��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�j(h�� ���Y�������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�j,h�� ���	�������t0�@,��t)�M$�E�UQ�M���\$�E�$R�UQR����^]�  3�^]�  �����������U��Vh�j0h�� ����������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh�j4h�� ���Y�������t5�@4��t.�M(�E �UQ�M���$R�UQ�MR�UQ�MRQ����^]�$ 3�^]�$ ������U��QVh�j8h�� �����������t�@8���E�t�E�MPQ���U�^��]� ��^��]� ����������U��Vh�j<h�� ����������t�@<��t�M�UQR����^]� ����������U��Vh�j@h�� ���i�������t�@@��t�M�UQR����^]� 3�^]� ���U��Vh�jHh�� ���)�������t�@H��t�M�UQR����^]� 3�^]� ���U��Vh�jDh�� �����������t�@D��t�M�UQR����^]� 3�^]� ���U��QVh�jLh�� ����������t#�@L���E�t�E�EP�����$�U�^��]� ��^��]� �����U��Vh�jPh�� ���Y�������t�@P��t�M�UQR����^]� 3�^]� ���U��Vh�jTh�� ����������t �@T��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�jXh�� �����������t(�@X��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh�j\h�� ���y�������t(�@\��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��V��~ Wu h�jh�� �"�������t�@�ЉF�~��t6h�jh�� ���������t�@��t�M�UVQ�MRQ����_^]� _3�^]� ��������������U��V��W�~��t+h�jh�� ��������t�@��t�M�UQR���Ѓ~ t1h�jh�� �p�������t�N�U�M�@R�Ѓ��F    _^]� ����������U��V��~ u h�jh�� �#�������t�@�ЉF�v��t+h�jh�� ���������t�@��t�M�UQR����^]� �������������U��V�q��t@h�jh�� ��������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ��������������U��V�q��t<h�j h�� �T�������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U��SV��~ Wu h�jh�� ��������t�@�ЉF�}�]�M�UWSQR���+  ��t�N��t�E�UWSPR����_^[]� _^3�[]� �U��V�q��t8h�j(h�� ��������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� ������U��I��t)�E$�E�UP�E���\$�E�$R�UPR����]�  3�]�  �������U��V�q��t<h�j0h�� ��������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U��E��u�E�M�����   ]� �����������U��E�����V��   �$����   ^]á�������uT�EP�#j����=�.  }�����^]Ëu��t�hP�jmh�j���������t ���iZ������tV���x^���   ^]���    �   ^]ËM�UQR�]������������^]�^]��c���-�u.��\����-������t����Z��V谹������    �   ^]Ã��^]Ð��?�F�����"�������������h�Ph�f �`������������������U��h�jh�f �<�������t
�@��t]�����]�������U��Vh�jh�f ����������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R��Y���E�NP�у�4�M����Y����^]ÍM��Y�����^]��U��h�jh�f ��������t
�@��t]��3�]��������U��h�jh�f �l�������t�x t�P]��3�]������V��F��Wu�~��N�ɍ<u�< ��u_3�^á`�H�F��  h��j8��    RP�у���tщ~�F_�   ^���U��V��F;Fu������u^]� �N�V�E���   F^]� �����������U��V��FW�};�~ ��|�F�M��_�   ^]� _3�^]� })�V;Vu��������t�F�N��    �F9~|׋V;Vu���������t��F�N�U���F_�   ^]� ������U��V��FW�};�~����}3�;Fu������u_^]� �F;�~�N�T������;ǉ�F�M���F_�   ^]� �U��E��|4�Q;�}-���;Q}V�d$ �Q�t������2;A|�^�   ]� 3�]� ������������U��Q3���V~�I�u91t����;�|���^]� �������V��W�~W����3����_�F�F^�����A    ��������̋Q�B���|;�}�QV�4���tP�1�����^�3�����������̍Q3��Q�Q�A�Q�A������������W���O�G;�t#��tV�q��t�~ u3���j�҅���u�^�G�G�G�G    �G�G    _�����U��A��3�;�Vt!��t�M���;�t�@��t
�x t��u�3�^]� ��������U��Q�E�P�Q�P�Q�B�A]� �U��E�Q�P�Q�P�Q�B�A]� ̋Q��3�;�t�ʅ�t�I����t
�y t��u�����������U��E�P�Q�H�A�@�H]� ����U��E�P�Q�H�A�A�H]� ���̋Q��t!�A��t�B�A�Q�P�A    �A    ��������V��W�~W�������3����_�F�F^��������������U���SV�uW���^S�}��ư��3���F�F�O�N�W���V9G�E~��I �O���F9F�U�uL��u�~��~��t���< ��t\�`�H���  h��j8��    RP�у���t3�~�}���V��M����E�F��;G�E|�_^�   [��]� _^3�[��]� �������������U��V�u��|'�A;�} �U��|;�};�t�A��W�<��<���_^]� ���������U��EV�u;�}����|,�Q;�}%��|!;�};�t�QW�<�P������tVW����_^]� ����������U��V�q3���W~�Q�}9:t����;�|���P�����_^]� ���������������U����E�Qj�E��ARP�M��E����|����]� �����U����Q�Ej�E��A�MRPQ�M��E�����|����]� ̋A��;�t?W3�;�t7V�H;�t	9yt���3��P;�t;�t�J�H�P�Q�x�x;���u�^_������̋Q�����t!�A��t�B�A�Q�P�A    �A    �̋�� ���@���HV3��q�q�P�r�r����p�p�p�P�H^������V����������F3�;��F��t�N;�t�H�F�N�H�V�V�F;��F��t�N;�t�H�F�N�H�V�V^�U��E�UP�AR�Ѓ�]� ���������U��V��N3�;����t�F;�t�A�F�N�H�V�V�Et	V薰������^]� ������������U��V��W�~W���*���3����E��F�Ft	V�Q�����_��^]� ������U��V��������Et	V�)�������^]� ���������������U��`�PH�EPQ���  �у�]� �U��`�P�B4VW�}j��h�  ���ЋMWQ���D  _^]� ��������������U��V���PXW�ҋ}P���������Et�_�   ^]� �M�UPWQR���1  _^]� �����������U��S�]VW��j �������8�  �}uI�~ uC�`�P���   j h�  ���Ѕ�u�`�QP���   h�  ���Ѕ�t	_^3�[]� �M�U�EQ�MRPSWQ����  _^[]� ��������U��EP�A    ��I����]� �����̸   �A� ������A   � ������U���@S�]��`��VW��u�G   �}  ����   �M3�V������8�  u4��@��P�w�I���`�P�M�B4��jh�  ��_^�C�[��]� �MV赸���8�  u�E�M��RPQ����_^�   [��]� �MV腸���8�  t�MV�t����8��  �`�P�M�B4jh�  �Љw�  ����  �E�H��BXj	��P�����3��؃�;މu�t�`�QH���  VS�Ѓ��E��M�;O�f  9w�]  �`�B�M���   Vh�  �҅�u!�`�P�M���   Vh�  �Ѕ��  �`�Q�M�B4Vh�  ��;�t
V���������E��G�`���   ���   �Ћ];މE���   ;���   S�'G���M���jQ�ˉu��uĉuȉủuЉu؉u���,���U�E��ˉu��u�u�U�E��]��E�   ��;����t!��t��t�u���E�   ��E�   ��E�   �a���M�;�t�>@����BX�M�Q����P�b���M܃�;�t�<@���M���v���M���v���M��H���]�M�U�EQSRP����  _^[��]� �M���G��_^�   [��]� �������������̸   � ��������� ������������̃��� ����������� �������������U��`�H�QV�uV�҃���^]� ̸   � ��������3�� ����������̸   @� ��������3��  ����������̸   � ��������U��W�}��u3�_]� ��U�@@VR�Ћ���u^_]� �`�Q0�F�M���   PQW�ҋF��^_]� U��`�H0�U�AR�Ѓ���t
��ȋj��]� �������3�� ��������������������������̸   � ��������3�� �����������3�� �����������U��E� ����]� �������������̸   � ��������U��E� ����]� ��������������3�� �����������U��`�H���  ]��������������U��`�H���  ]��������������U��`�P�EP�EP�EP�EPQ���   �у�]� �����U��`�E�P�EP�E���\$�E�$PQ���   �у�]� �������������U��`�P�EP�EP�EPQ���   �у�]� ��������̡`�P���   Q�Ѓ�������������U��`�P�EP�EP�EPQ���   �у�]� ���������U��`�P�EP�EPQ���   �у�]� �������������U��`�H�U�ApR�Ѓ�]� �����U��`�P�EP�EPQ���  �у�]� �������������U��`�P�EP�EPQ���  �у�]� �������������U��`�P�EP�EPQ���  �у�]� �������������U��`�P�EP�EPQ���  �у�]� �������������U����   V�u��u3�^��]�Wh�   ��0���j P��  ��R���E�P���ҡ`�P�B<�M��Ѕ��}t0j �M�QW��������u�`�B�P�M�Q�҃�_3�^��]ËE�M�Uh�   ��p�����0���P��t����MQWj	��P�����0���ǅ4���k �E���E�@��E����E� �E���E���E�p�ǅx����o ǅ|����o �E���E��E���E�P��E����E� ��E� ��E�`��E� �E�0��E��o ��Z���`���B�P�M�Q�҃�_��^��]����������U���   SV�u(3ۅ��]�u�`�H�A�UR�Ѓ�^3�[��]Ë`�Q�B<W�M3��Ѕ��'  謓�����E�tq�MQ�M��YF��Wh���M��B��P�M��BF���u�Wj��U�R�E�P��\���Q�_?�eX����P��x���R��I����P�E�P��I����P���������E�t�E� �� t�M�����`F����t��x�������MF����t��\�������:F����t�M̃���*F����t�`�Q�J�E�P����у���t�M�� F���}� t"�U(�E$�M�R�UP�EQ�MRPQ���������U�R蟒������E$�M�UVP�Ej QRP����������`�Q�J�EP�у���_^[��]����������������U��E�M�UP�EQ�Mj RPQ������]�������������̋�`L����������̋�`0����������̋�`P����������̋�`����������̋�`$����������̋�`D����������̋�`T����������̋�`����������̋�`(����������̋�`HQ���a  Y�V��������D$tV�h���Y��^� U��Q�E��SVW�  ����   Wj ��P������u3��  V�>����Vj u��P���ދF�~�E�F�E�F�E����  ��P���E��t�� �  �M����E�����j�������=��-  ��Y�s����$  ��u
�p  �`����i  ����$�$  ���N  ��}��  ���Q  ��| ��  ��|j �R  ��Yu���   �i  ��3�;�u59=��������9=	u�  9}u{�8  �s  ��  �j��uY�0  h  j�/  ��;�YY�����V�5$��5 	�  Y�Ѕ�tWV�g  YY� ��N���V�  Y�m�����uW�  Y3�@_^[�� jh@��D   ����]3�@�E��u9���   �e� ;�t��u.����tWVS�ЉE�}� ��   WVS������E����   WVS�L����E��u$��u WPS�8���Wj S��������tWj S�Ѕ�t��u&WVS�~�����u!E�}� t����tWVS�ЉE��E������E���E��	PQ�T  YYËe��E�����3��  Ã|$u�L!  �t$�L$�T$�����Y� �U � ���Q������C���������������� �9��$����������-  �|$ ��t�k-  ���;��u����-  ���̃=�# t-U�������$�,$�Ã=�# t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$���5���  ��Yt��j�H/  jj �!/  ���&.  �����������U��WV�u�M�}�����;�v;���  ��   r�=�# tWV����;�^_u^_]�O1  ��   u������r*��$�����Ǻ   ��r����$����$�����$�(�������#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ���������r���$����I ��x�p�h�`�X�P�H��D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��������������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�0������$����I �Ǻ   ��r��+��$�4��$�0��D�h����F#шG��������r�����$�0��I �F#шG�F���G������r�����$�0���F#шG�F�G�F���G�������V�������$�0��I �����������'��D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�0���@�H�X�l��E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_������������̋T$�L$��ti3��D$��u��   r�=�# t�4/  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$�jh`���  �e� �u;5�#w"j��0  Y�e� V�9  Y�E��E������	   �E���  �j��/  Y�U�l$�����   S��VW3�95<
��u�k,  j��*  h�   ��  YY��#��u;�t���3�@P���uU�S���;�Yu;�u3�G�����WV�5<
�Ӌ���u&9�j_tU��;  ��Yu���j;  �8�c;  �8_��^[]�U�;  Y�N;  �    3�]�jh����  �u��tu�=�#uCj�/  Y�e� V�$0  Y�E��t	VP�@0  YY�E������   �}� u7�u�
j�.  Y�Vj �5<
����u��:  ����P�:  �Y�  ������̃=�# ��=  ���\$�D$%�  =�  u�<$f�$f��f���d$��=  � �~D$f(0�f(�f(�fs�4f~�fT`�f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�f:  ���D$��~D$f��f(�f��=�  |!=2  �fT ��\�f�L$�D$����f�P�fVP�fT@�f�\$�D$�QSUVW�5�$�  �5�$���t$��  ��;�YY��   ��+ލk��rxV�A=  ��;�YsJ�   ;�s���;�rP�t$�  ��YYu�F;�rCP�t$�h  ��YYt3��P�<��  Y��$�t$�  ���W��  Y��$�D$Y�3�_^][Y�Vjj ��  ��V��  ������$��$ujX^Ã& 3�^�jh���#  �  �e� �u�����Y�E��E������	   �E��?  ��|  ��t$���������YH���������̃��$�?  �   ��ÍT$�H?  R��<$�D$tQf�<$t� ?  �   �u���=� �s?  �   ����p?  �  �u,��� u%�|$ u����>  �"��� u�|$ u�%   �t����-���   �=� �?  �   ����>  Z������̺���a@  �����?  �Ƀ=�t����TL  �����z����jh����  j��+  Y�e� �u�N��t/�����E��t9u,�H�JP�����Y�v�����Y�f �E������
   ��  Ë���j�*  Y��������������̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t������&  �t$�6%  �5 ���  h�   �Ѓ��h��� ���thp�P����t�t$����t$�����Y�t$�$��j�*  Y�j�)  Y�V������t�Ѓ�;t$r�^�V�t$3����u���t�у�;t$r�^ËL$V3�;�u�5  VVVVV�    � O  ��jX^á�;�tډ3�^ËD$V3�;�u�h5  VVVVV�    ��N  ��jX^�95�tۋ��3�^Ã=� th��9P  ��Yt�t$��Y�*!  hD�h,��6�����YYuTVWh!������ ��ƿ(�;�Ys���t�Ѓ�;�r�=�$ _^th�$��O  ��Ytj jj ��$3��jh���&  j�,)  Y3��}�3�C9	t~�	�E�	9}u[�5�$��  �E��5�$��  YY���u�9}�t&���u�;u�r�> t��>�  ;�t�W�  Y����hT��H��2���Yh\��X��"���Y�E������   �} u(�	j�'  Y�u�����3�C�} tj�'  Y��  �j j�t$�������jj j �������V�   ��V��3  V�Q  V��K  V�M$  V�Q  V�O  V�  V�tO  h���v   ��$� �^�U��QQSV3��E�F3�P�u��]�������}�Y~���BWS� ��p<�f9^�F�|0v#Wh���0�����YYt�FC��(;�r���e� �E�_^[��V�5(��5(��օ�t!�$����tP�5(����Ѕ�t���  �&h��� �����t#�J�����th��V����t
�t$�ЉD$�D$^�j ����Y�V�5(��5(��օ�t!�$����tP�5(����Ѕ�t���  �&h��� �����t#�������th��V����t
�t$�ЉD$�D$^��,�� V�5(��(�����u�5	�k���Y��V�5(��0���^á$����tP�5$	�A���Y�Ѓ$���(����tP�4��(����$  jh ��  h��� ��E�u�F\x�3�G�~��t/������t&h���u���Ӊ��  h���u��Ӊ��  �~pƆ�   CƆK  C���FhP�8�j�%  Y�e� �E�Fl��u����Fl�vl�8Q  Y�E������   �  �j�$  Y�VW���5$��������Ћ���uNh  j�  ����YYt:V�5$��5 	����Y�Ѕ�tj V�����YY� ��N���	V�(���Y3�W�<�_��^�V��������uj�����Y��^�jh ���  �u����   �F$��tP�����Y�F,��tP�����Y�F4��tP�����Y�F<��tP����Y�FD��tP����Y�FH��tP����Y�F\=x�tP����Yj�W$  Y�e� �~h��tW�@���u���tW�Y���Y�E������W   j�$  Y�E�   �~l��t#W�BP  Y;=��t�� �t�? uW�`N  Y�E������   V����Y�  � �uj��"  YËuj��"  YÃ=$��tLW�|$��u&V�5(��5(��օ�t�5$��5(����Ћ�^j �5$��5 	�`���Y��W����_�(����t	j P�0��Wh��� �����u	�����3�_�V�5�h�W��hظW�	��h̸W�	��hĸW� 	�փ=	 �50��$	t�=	 t�= 	 t��u$�(��	�4��	U��5 	�$	�,�����(���   �5	P�օ���   �J����5	������5	�	������5 	�	������5$	� 	��������$	��   ��teh��5	����Y�Ѓ���$�tHh  j�   ����YYt4V�5$��5 	�����Y�Ѕ�tj V�����YY� ��N��3�@��l���3�^_�VW3��t$�#�������Yu'9(	vV�D����  ;(	v��������uɋ�_^�VW3�j �t$�t$�U  ������u'9(	vV�D����  ;(	v��������u���_^�VW3��t$�t$�V  ����YYu-9D$t'9(	vV�D����  ;(	v��������u���_^�jThH���	  3��}��E�P�T��E�����j@j ^V�@���YY;��  ��#�5�#��   �0�@ ���@
�x�@$ �@%
�@&
�x8�@4 ��@��#��   ;�r�f9}��
  �E�;���   �8�X�;�E�   ;�|���E�   �[j@j ����YY��tV�M����#���# ��   �*�@ ���@
�` �`$��@%
�@&
�`8 �@4 ��@��;�r��E�9=�#|���=�#�e� ��~m�E����tV���tQ��tK�uQ�P���t<�u���������4��#�E� ���Fh�  �FP�/I  YY����   �F�E�C�E�9}�|�3ۋ���5�#����t���t�N��r�F���uj�X�
��H������P�L������tC��t?W�P���t4�>%�   ��u�N@�	��u�Nh�  �FP�H  YY��t7�F�
�N@�����C���g����5�#�H�3��3�@Ëe��E����������  �VW��#�>��t1��   �� t
�GP�X����@   ;�r��6�����& Y�����$|�_^�S3�9�$VWu�_R  �5�3�;�u����   <=tGV�C  Y�t�:�u�jGW������;�YY�=�tˋ5�U�@V�bC  ��E�>=Yt/jU�Z���;�YY�tJVUP��B  ����tSSSSS�A  �����8u��5�����������$   3�Y]_^[��5������������U��Q�MS3�9EV���U�   t	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF��T  ��Yt��} t
�M��E�F�ۋU�Mt2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=����Pt#�T  ��Yt��M�E�F��M��E����S  ��YtF���UF�V�����t� B�U��M�����E��^[t�  ���U���S3�9�$VWu��O  h  �0	VS�4
�\���$;É5	t8�E�u�u��U��E�PSS�}������E���=���?sJ�M���sB�����;�r6P������;�Yt)�U��E�P�WV�}�������E���H���5�3�����_^[��QQ�8
SUVW�=p�3�3�;�j]u-�׋�;�t�8
   �"����xu	�ţ8
��8
����   ;�u�׋�;�u3���   f9��t�f9u��f9u�=l�SSS+�S��@PVSS�D$4�׋�;�t2U�����;�Y�D$t#SSUP�t$$VSS�ׅ�u�t$����Y�\$�\$V�h����X;�t;�u��d���;��p���8t
@8u�@8u�+�@��U�Z�����;�YuV�`��D���UVW�6�����V�`���_^][YY�VW�0��0�;ǋ�s���t�Ѓ�;�r�_^�VW�8��8�;ǋ�s���t�Ѓ�;�r�_^�U��QQV�E�3�P�u��u��U�����YtVVVVV�j=  ���E�P�q�����YtVVVVV�O=  ���}�^u�}�r3�@��jX��3�9D$j ��h   P�x����<
u3���}�������#u$h�  �J  ��Yu�5<
�t��%<
 ��3�@�U3�=�#uTS��W3�9-�#~1V�5�#��h �  U�v��|��6U�5<
�Ӄ�G;=�#|�^�5�#U�5<
��_[�5<
�t��-<
]��U��QQV���������F  �V\���W�}��S99t��k����;�r�k��;�s99u���3���t
�X�ۉ]�u3���   ��u�` 3�@��   ����   �N`�M��M�N`�H����   ����=�����;�}$k��~\�d9 �=�����B߃�;�|�]�� =�  ��~du	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=�  �u	�Fd�   �=�  �u�Fd�   �vdj��Y�~d��` Q�ӋE�Y�F`���[_^�øcsm�9D$u�t$P����YY�3��hP�d�5    �D$�l$�l$+�SVW���1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q���������������̃�S�\$ UV�s35��W�����D$ �D$   �{t�N�38�����N�F�38�����D$(�@f�  �k����L$0�T$�D$�L$ �S�t^�Dm �L��ɍ\���D$t����N  ���D$|DL�D$�����ù|$ t$����t�N�38�����N�F�38�����D$_^][����D$    �ƋL$(�9csm�u*�=�# t!h�#�<  ����t�T$(jR��#���L$,�vN  �D$,9hth��W�Ջ��xN  �D$,�L$�H����t�N�38�����N�V�3:�r����K���N  �{��P���h��W�˺�����#N  ����U�������e� �e� SW�N�@�;ǻ  ��t��t	�У���`V�E�P����u�3u����3�� �3����3��E�P����E�3E�3�;�u�O�@����u������5���։5��^_[��U��� S3�9]u ��  SSSSS�    �49  ������   �M;�V�ut!;�u�  SSSSS�    �9  ������S����;ȉE�w�M�W�u�E��u�E�B   �u�u�P�u��O  ��;��t�M�x�E����E�PS��L  YY��_^[���t$j �t$�t$�t$�8�����ËD$��V���F uc�����F�Hl��Hh�N�;��t�0��Hpu�v@  ��F;0�t�F�0��Hpu��B  �F�F�@pu�Hp�F�
���@�F��^� U���V�u�M��l����u�P�Y  ��e�F�P�7X  ��Yu��P�iY  ��xYuFF�M����   �	��	�F�����F��u�8M�^t�E��`p���U���V�u�M�������E��ɋu�t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B�Ɉu��}� ^t�E��`p�����D$�����Az3�@�3��U��QQ�} �u�ut�E�P�X  �M��E��M��H��EP�7Y  �E�M�����j �t$�t$�t$������Å�V��tV�-7  @PV�V�Y  ��^�j �t$�z���YY�j �t$�����YY�U���SVW�u�M��������3�;�u+��  j_VVVVV�8�B6  ���}� t�E��`p����!  9uv�9u~�E�3���	9Ew	�  j"뺀} t�U3�9u��3Ƀ:-����ˋ��:����}�?-��u�-�s�} ~�F�����E����   � � �3�8E��E��}�u����+�]h�SV�5  ��3ۅ�tSSSSS�4  ��9]�Nt�E�GF�80t.�GHy���-F��d|
�jd_�� ��F��
|
�j
_�� �� F��t�90uj�APQ�+X  ���}� t�E��`p�3�_^[��U���,���3ŉE��ESVW�}j^V�M�Q�M�Q�p�0��\  3ۃ�;�u�W  SSSSS�0�4  �����o�E;�v����uu����3Ƀ}�-��+�3�;���+��M�Q�NQP3��}�-��3�;�����Q��Z  ��;�t���u�E�SP�u��V�u��������M�_^3�[������U��j �u�u�u�u�u������]�U���$VW�u�M��E��  3��E�0   �k���9}}�}�u;�u+�q  j^WWWWW�0��3  ���}� t�E�`p����  9}vЋE��9E� w	�3  j"���}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW� �������t�}� � ��  �M�ap��  �;-u�-F�0F�} je����$�x�FV��R  ��YY�L  �} ���ɀ����p��@ �2  %   �3��t�-F�]�0F������$�x��OF��ۃ����  �3���'3��u!�0�O����� F�u�U���E��  ��1F��F9U�Eu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~M�W#U���M�#E���� �[  f0 ��f=9 vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �5[  f= v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V�M�����u�E�8 u���} �4����$�p���WF��Z  3�%�  #�+E�SY�x;�r�+F�
�-F�����;Ӌ��0|$��  ;�rSQRP�Y  0�F;��U�����u��|��drj jdRP�vY  0��U�F����;�u��|��
rj j
RP�PY  0��U�F���]�0��F �}� t�E�`p�3�[_^��U���SVW�u�؋s���M�N������u-�  j^�03�PPPPP�r0  ���}� t�E��`p����   �} v̀} t;uu3��;-����� 0�@ �;-��u�-�w�C3�G�����n����0F���} ~D���Y����E����   � � ��[F��}&�ۀ} u9]|�]�}���(���Wj0V�������}� t�E��`p�3�_^[��U���,���3ŉE��ESVW�}j^V�M�Q�M�Q�p�0�pW  3ۃ�;�u�  SSSSS�0�j/  �����Z�E;�v���u��3Ƀ}�-��+��u�M�Q�M��QP3��}�-���P�U  ��;�t���u�E�SV�u���d������M�_^3�[�X�����U���0���3ŉE��ESV�uWj_W�M�Q�M�Q�p�0�V  3ۃ�;�u�L  SSSSS�8�.  �����   �M;�vދE�H�E�3��}�-������<0u��+ȍE�P�uQW��T  ��;�t��X�E�H9E������|-;E}(:�t
�G��u��_��u�E�j�u���u��������u�E�jP�u���u�u�������M�_^3�[�`�����U��E��et_��EtZ��fu�u �u�u�u�u�&�����]Ã�at��At�u �u�u�u�u�u�����0�u �u�u�u�u�u������u �u�u�u�u�u�|�����]�U��j �u�u�u�u�u�u�^�����]�VW3��� ��6���������(Y�r�_^�Vh   h   3�V�V  ����tVVVVV�,  ��^�U���� ��]�����]��E��u��M��m��]����]�����z3�@��3���h$�� ���th�P����tj �������U���(  �H�D�@�<�58�=4f�`f�Tf�0f�,f�%(f�-$��X�E �L�E�P�E�\��������
  �P�L
�@
	 ��D
   �����������������������
j��U  Yj ���h0�����=�
 uj�U  Yh	 ����P����Ã%�# ��U  ��#3��U��$X�����(  ���3ŉ��  �(�Vtj
��   Y�U.  ��tj�W.  Y�(���   ���   ���   ���   �]|�ux�}tf���   f���   f�]pf�Elf�ehf�md����   ���  ���  ���   �E�  ���   �@�jP���   �E�j P�����E����EЍE�j �E�  @�u��E�����E�P���j�k���̋L$�(��T$#T$��#�ʉ(��QS�\$VW3�3�;�0�tG��r���w  Uj��W  ��Y�1  j��W  ��Yu�=��  ���   �?  h��  S�hU�8*  ����tVVVVV�)  ��h  ��Vj �� �\���u&hȾh�  V��)  ����t3�PPPPP��(  ��V�E*  @��<Yv8V�8*  ��;�j�|hľ+�QP�sV  ����t3�VVVVV�(  ���3�h��SU��U  ����tVVVVV�\(  ���4�4�SU�U  ����tVVVVV�:(  ��h  h��U��S  ���3j��L���;�t%���t j �D$P�4�4��6�)  YP�6U���]_^[Y�j�uV  ��Ytj�hV  ��Yu�=�uh�   �4���h�   �*���YYËD$���U����}��u��u�}�M�����    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Iu��u��}���]�U����}�u��]��]�Ù�ȋE3�+ʃ�3�+ʙ��3�+���3�+����uJ�u�΃��M�;�t+�VSP�'������E�M��tw�]�U�+щU��+ى]��u�}��M��E�S;�u5�ك��M�u�}�M��MM�UU�E+E�PRQ�L������E��u�}�M�����ʃ��E�]��u��}��]�U����}��}�M��f�����$    �ffGfG fG0fG@fGPfG`fGp���   IuЋ}���]�U����}��E���3�+���3�+���u<�M�у��U�;�t+�QP�s������E�U��tEE+E�3��}��M��E�.�߃��}�3��}�M��E��M�U�+�Rj Q�~������E�}���]�VW3����<���u�����8h�  �0����*  ��YYtF��$|�3�@_^Ã$��� 3���S�X�V���W�>��t�~tW��W�1����& Y�����|ܾ��_���t	�~uP�Ӄ����|�^[�U��E�4������]�jhh�����3�G�}�3�9<
u����j�����h�   �����YY�u�4���9t���nj����Y��;�u��  �    3��Qj
�Y   Y�]�9u,h�  W��)  YY��uW�a���Y�  �    �]���>�W�F���Y�E������	   �E��B����j
�*���Y�U��EV�4����> uP�$�����Yuj�����Y�6���^]�h@  j �5<
������#uËL$�%� �%�# ��#3���#��#   @Ë�#��#k����T$+P��   r	��;�r�3��U����M�AV�uW��+y�������i�  ��D  �M��I���M���  S�1��U�V��U��U����]ut��J��?vj?Z�K;KuB�� �   �s����L��!\�D�	u#�M!��J���L��!���   �	u�M!Y�]�S�[�M�M�Z�U�Z�R�S�M�����J��?vj?Z�]����]���   +u��]���j?�uK^;�v��M�����J;։M�v��;�t^�M�q;qu;�� �   �s������!t�D�Lu!�M!1��K�����!���   �Lu�M!q�M�q�I�N�M�q�I�N�u��]�}� u;���   �M��ыY�N�^�q�N�q�N;Nu`�L�M���� �Ls%�} u�ʻ   ���M	�   �����D�D	�)�} u�J�   ���M	Y�J�   ��ꍄ��   	�E���D0��E����   ������   ��#�5|�h @  ��H� �  SQ�֋�#���   ���	P���@��#����    ���@�HC���H�yC u	�`����x�ueSj �p�֡��pj �5<
����#��k���#+ȍL�Q�HQP�hD  �E����#;�v�m��#��#�E���=�#[_^�á�#V�5�#W3�;�u4��k�P�5�#W�5<
���;�u3��x��#�5�#��#k�5�#h�A  j�5<
��;ǉFt�jh    h   W���;ǉFu�vW�5<
��뛃N��>�~��#�F����_^�U��QQ�M�ASV�qW3���C��}���i�  ��0D  j?�E�Z�@�@��Ju�j��h   ��yh �  W�����u����   �� p  ;��U�wC��+����GA�H�����  ����  ��������@��  �Pǀ�  �     IuˋU��E��  �O�H�A�J�H�A�d�D 3�G����   �FC�������E�NCu	x�   �������!P��_^[��U����M�ASV�uW�}��+Q������i�  ��D  �M�O����I;�|9���M�]��U  ���E  �;��;  �M���I��?�M�vj?Y�M��_;_uC�� �   �s��M��L��!\�D�	u&�M!������M��L��!���   �	u�M!Y�O�_�Y�O��y�M+�M��}� ��   �}��M��O��?�L1�vj?_�]���]�[�Y�]�Y�K�Y�K�Y;YuW�L�M���� �Ls�} u�ϻ   ���M	�D�D��� �} u�O�   ���M	Y����   �O�   ���	�U�M��D2���L���U�F�B��D2��<  3��8  �/  �])u�N�K��\3��u��N��?�]�K�vj?^�E���   �u���N��?vj?^�O;OuB�� �   �s����t��!\�D�u#�M!��N���L��!���   �	u�M!Y�]�O�w�q�w�O�q�uu��u��N��?vj?^�M��y�K�{�Y�K�Y�K;KuW�L�M���� �Ls�} u�ο   ���M	9�D�D��� �} u�N�   ���M	y����   �N�   ���	�E��D�3�@_^[��U�����#�Mk��#������M���SI�� VW}�����M���������3���U���#����S�;#U�#��u
��;؉]r�;�u��#��S�;#U�#��u
��;ى]r�;�u[��{ u
���];�r�;�u1��#�	�{ u
��;ى]r�;�u�����؅ۉ]u3��	  S�@���Y�K��C�8�t��#�C�����U�t����   �|�D#M�#��u)�e� ���   �HD�9#U�#��u�E����   ����U���i�  ��D  �M�L�D3�#�u����   #M�j _��G��}��M�T��
+M�����N��?�M�~j?^;��  �J;Ju\�� �   �}&����M��|8�Ӊ]�#\�D�\�D�u3�M�]!�,�O���M�����   �|8��!��]�u�]�M�!K��]�}� �J�z�y�J�z�y��   �M��y�J�z�Q�J�Q�J;Ju^�L�M���� �L}#�} u�   �����	;�ο   ���M�	|�D�)�} u�N�   ���	{�M�����   �N�   ���	7�M���t�
�L���M��u�эN�
�L2��u��ɍy�>u;�u�M�;�#u�%� �M���B_^[�ËD$3�;��tA��-r�H��wjXË���D���jY;��#�����'�����u�p�Ã��������u�t�Ã��V������L$Q�����Y��������0^ËD$����5��.�����Yt�t$�Ѕ�Yt3�@�3��U���(3�9�S�]V�uW�}�E��E��E��E��E��E��E��E�t�5�#�����Y���[�M��   ;��t  �[  ����   ��   ��jY+���   J��   ����   J��   ��tqJtE��	��  �E�   �Eܼ���M��]�Q��]���]��Ѕ�Y��  ����� "   �  �Eܸ���M��]�Q��E�   �]���]���Y�j  �E�   �Eܸ���Eܰ���]���]���"  �M��Eܰ��r����Eܬ��׉M��Eܬ��Z����Eܼ�놃�tNIt?It0It ��t����   �Eܤ���Eܜ���Eܼ�����Eܼ��x����E�   ��������   �E�   �Eܔ���������������   �$�L�Eܬ���Eܰ���Eܸ���E܌���E܄���E�|��y����E�t��m����E�p���E�l���E�h���M����]���]�M��]�Q�E�   �Ѕ�Yu�&���� !   �E��_^[�Ë�������i�SJ��U��QQSV���  V�5x��lL  �EYY�؋EQf%�f=�Q�$uU�-K  ��YY~-��~��u#�ESQQ�$j��I  ���rVS�"L  �EYY�d�ES�����\$�E�$jj�?�J  �]��EY�]�Y����DzVS��K  �E�YY�"�� u��E�S���\$�E�$jj�I  ��^[��jh������3��]3�;���;�u������    WWWWW�O  ������S�=�#u8j�[���Y�}�S�����Y�E�;�t�s���	�u���u��E������%   9}�uSW�5<
��������K����3��]�u�j�+���Y������������̀zuf��\���������?�f�?f��^���٭^�������剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^�������剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp���������۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-����p��� ƅp���
��
�t���������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR��I  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   �����   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z��������������ܿ�����   s������������������Կ�����   v���������U���0���S�ٽ\�����=@� t������8����   [����ݕz������U���U���0���S�ٽ\����=@� t�������8�����8�����Z   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���ƅq���������   [�À�8�����=� uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   �(�����������������s4�8��,ǅr���   � �����������������v�0�VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�/F  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8������������[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[���l$�l$�D$���   5   �   t��������� u��ËD$%�  tg=�  t`�|$�D$?  %��  �D$ �l$ �D$%�  ��t�����������l$��������������l$��ËD$D$u��ËD$%�  u��|$�D$?  %��  �D$ �l$ �D$%�  t=�  t2�D$�s*��D$�r ����������|$�l$�ɛ�l$������l$��Ã�,��?�$������,Ã�,�����,Ã�,�����,�����,�����,�����,��|$���<$�|$ �����l$ �Ƀ�,Ã�,��<$�|$�����l$�Ƀ�,Ã�,����|$���<$�|$ �^����l$ ��,��<$�|$�J�����,��|$�<$�:����l$��,��|$�<$�&�����,��|$�����<$�|$ �������l$ �ʃ�,Ã�,��<$���|$��������l$�ʃ�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$�����Ƀ�,��|$���<$�������l$��,��|$���<$�����Ƀ�,��|$�����<$�|$ �j������l$ �˃�,Ã�,��<$���|$�K������l$�˃�,Ã�,����|$�����<$�|$ �$������l$ ��,��<$���|$�����ʃ�,��|$���<$��������l$��,��|$���<$������ʃ�,��|$�����<$�|$ ��������l$ �̃�,Ã�,��<$���|$�������l$�̃�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�h����˃�,��|$���<$�T������l$��,��|$���<$�<����˃�,��|$�����<$�|$ �"������l$ �̓�,Ã�,��<$���|$�������l$�̓�,Ã�,����|$�����<$�|$ ��������l$ ��,��<$���|$������̃�,��|$���<$�������l$��,��|$���<$�����̃�,��|$�����<$�|$ �~������l$ �΃�,Ã�,��<$���|$�_������l$�΃�,Ã�,����|$�����<$�|$ �8������l$ ��,��<$���|$� ����̓�,��|$���<$�������l$��,��|$���<$������̓�,��|$�����<$�|$ ��������l$ �σ�,Ã�,��<$���|$�������l$�σ�,Ã�,����|$�����<$�|$ �������l$ ��,��<$���|$�|����΃�,��|$���<$�h������l$��,��|$���<$�P����΃�,Ã�,�<$�|$�;�����,Ã�,�|$�<$�(�����,�P�D$%  �=  �t3��% 8  t�D$����X� �Ƀ��<$�D$�����,$�Ƀ�X� �t$X� P�D$%  �=  �t3��% 8  t�D$�k���X� �Ƀ��<$�D$�V����,$�Ƀ�X� �t$X� P��% 8  t�D$�/���X� �Ƀ��<$�D$�����,$�Ƀ�X� P��% 8  t�D$�����X� �Ƀ��<$�D$������,$�Ƀ�X� P�D$%  �=  �t3��% 8  t�D$�����X� �Ƀ��<$�D$�����,$�Ƀ�X� �|$X� P�D$%  �=  �t3��% 8  t�D$�~���X� �Ƀ��<$�D$�i����,$�Ƀ�X� �|$X� P��% 8  t�D$�B���X� �Ƀ��<$�D$�-����,$�Ƀ�X� P��% 8  t�D$����X� �Ƀ��<$�D$������,$�Ƀ�X� P��,�<$�|$������,X�P��,�|$�<$�������,X�PSQ�D$5   �   ��  �������� �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u��������Ƀ�u�\$0�|$(���l$�-������l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8����l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$3ҋD$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w������|$����<$� �|$$�D$$   �D$(�l$(������<$�l$$�T�����0Z�����0Z�PSQ�D$5   �   ��  �������� �p  �D$%  �=  ��\  �D$.%  ��M  =  ��B  �D$,��6  �D$��*  �D$%�  ��?�\$0���  +�w^�D$%�  ��
�\$0���  +���   �l$(�D$�\$0���  ��+؃���+ˋ؁� �  ˉL$�l$�D$�����|$(�����   u�l$�|$�|$4�D$4?  �D$8�l$8�D$%�  �\$0���  +؃�?�� ���ˋD$�\$0���  % �  ؉\$�l$���l$(������%   u��������Ƀ�u�\$0�|$(���l$�-������l$(�l$4�� �  t���
�l$�l$(����   tV�|$<��   t�|$4�D$4   �D$8�l$8����l$4�D$<�����l$��% C  ���4$�d$��  	D$�$$��Y[X�R��0�|$�<$�    �D$�  �t
�������0Z��,$�l$�$D$ty���|$�,$�Ƀ��|$$�D$$?  �D$(�l$(�D$ %�  =�  w������|$����<$� �|$$�D$$   �D$(�l$(������<$�l$$�Q�����0Z�����0Z�������@���������ËD$���U��$X�����(  ���3ŉ��  V���   ���   ���   �]|�ux�}tf���   f���   f�]pf�Elf�ehf�md����   ���  ���  ���   �E�  ���   �@�jP���   �E�j P�*����E��EЍE؃��E�  ��u��E����j ������E�P�����u��uj�*  Yh  ����P������  3�^�d����Ũ  ��U���5�������Yt]��j��)  Y]������L$S3�;�VWt�|$;�w�Q���j^�0SSSSS���������1�t$;�u��ًъ�BF:�tOu�;�u�����j"Y�����3�_^[������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+������̋L$f�9MZt3�ËA<��8PE  u�3�f�x�����������̋D$�H<��ASV�q3҅�W�Dv�|$�H;�r	�X�;�r����(;�r�3�_^[���������������U��j�h��hP�d�    P��SVW���1E�3�P�E�d�    �e��E�    h   �<�������tU�E-   Ph   �R�������t;�@$���Ѓ��E������M�d�    Y_^[��]ËE��3�=  ���Ëe��E�����3��M�d�    Y_^[��]�jh�������ǳ���@x��t�e� ���3�@Ëe��E����������������h+0����Y�(ËD$�,�0�4�8ËD$���V9Pt��k�t$��;�r�k�L$^;�s9Pt3���54����Y�j h������3��}�}؋]��Lt��jY+�t"+�t+�td+�uD腲�����}؅�u����a  �,�,�`�w\���`���������Z�Ã�t<��t+Ht�����    3�PPPPP�t�����뮾4�4��0�0�
�8�8�E�   P�V����E�Y3��}���   9E�uj����9E�tP�=���Y3��E���t
��t��u�O`�MԉG`��u@�Od�M��Gd�   ��u.����M܋������9M�}�M�k��W\�D�E���辯����E������   ��u�wdS�U�Y��]�}؃}� tj �����Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3�诿��ËD$�@ËD$�D��t$���3�@� jh��9���3��}��5D�(���Y��;�uS�E�P����Y;�tWWWWW��������}�t!h��� �;�thX�P����;�u��2V�]���Y�D�}��u�u�։E��/�E� � �E�3�=  �����Ëe�}�  �uj�<��e� �E������E��ƾ���SUV�t$���   3�;�Wto=Hth���   ;�t^9(uZ���   ;�t9(uP�w������   ��4  YY���   ;�t9(uP�V������   �4  YY���   �>������   �3���YY���   ;�tD9(u@���   -�   P�������   ��   +�P��������   +�P�������   ���������   �=� t9��   uP�2  �7迤��YYj�~P[���t�;�t9(uP螤��Y9o�t�G;�t9(uP臤��Y��Ku�V�z���Y_^][�SUV�t$W�=8�V�׋��   ��tP�׋��   ��tP�׋��   ��tP�׋��   ��tP��j�^P]�{��t	���tP�׃{� t
�C��tP�׃�Mu؋��   �   P��_^][�V�t$��tSUW�=@�V�׋��   ��tP�׋��   ��tP�׋��   ��tP�׋��   ��tP��j�^P]�{��t	���tP�׃{� t
�C��tP�׃�Mu؋��   �   P��_][��^Å�t7��t3V�0;�t(W�8�������YtV�R����> Yu�� �tV�x���Y��^�3��jh(������������0��Fpt"�~l t�����pl��uj �ڧ��Y��������j����Y�e� �Fl�=���i����E��E������   ��j����Y�u��-�  t"��t��tHt3�ø  ø  ø  ø  �SUVW�  ��U3��^WS�۠���~�~�~3��~�������+Ɗ�CMu���  �   ��ANu�_^][�U��$d�����  ���3ŉ��  SW�E�P�v�İ���   ��   3����  @;�r�E���ƅ�   t+�]����;�w+�@P���  j R�+�����C�C��u�j �v�E��vPW���  Pjj �3  3�S�v���  WPW���  PW�vS�7  ��DS�v���  WPW���  Ph   �vS�7  ��$3��LE���t�L���  ���t�L ���  ��  �Ƅ   @;�r��M��  �E�����3�)E��U���  ЍZ ��w�L�р� ���w�L �р� ���  A;�rŋ��  _3�[蹚���Ŝ  ��jhH��`����v������0��Gpt�l t�wh��uj �[���Y���x����j�8���Y�e� �wh�u�;50�t6��tV�@���u���tV�/���Y�0��Gh�50��u�V�8��E������   뎋u�j�����Y�U���S3�S�M���������lu�l   �̰8]�tE�M��ap��<���u�l   �Ȱ�ۃ��u�E��@�l   ��8]�t�E��`p���[��U��� ���3ŉE�S�]V�uW�h�����3�;��}u�������3��  �u�3�9�8���   �E��0=�   r����  �f  ����  �Z  ��P�а���H  �E�PW�İ���)  h  �CVP�U���3�B��9U�{�s��   �}� ��   �u�����   �F����   h  �CVP�����M��k�0�u���H��u��*�F��t(�>����E���4�D;�FG;�v�}FF�> uыu��E����}��u�r�ǉ{�C   ����j�C�C��<�Zf�1Af�0A@@Ju������������L@;�v�FF�~� �4����C��   �@Iu��C�.����C�S��s3��{����95l�b�������M�_^3�[輗����jhh��i����M���{������}�������_h�u�����E;C�W  h   �v���Y�؅��F  ��   �wh���# S�u�����YY�E�����   �u��vh�@���u�Fh=�tP����Y�^hS�=8����Fp��   �0���   j�����Y�e� �C�|�C���C��3��E��}f�LCf�Ep@��3��E�=  }�L��(�@��3��E�=   }��  ��0�@���50��@���u�0�=�tP�`���Y�0�S���E������   �0j�B���Y��%���u ���tS�*���Y�h����    ��e� �E��!���Ã=�$ uj��V���Y��$   3��jh��豴���M3�;�v.j�X3���;E�@u�����    WWWWW�m�����3���   �M��u;�u3�F3ۉ]���wi�=�#uK������u�E;�#w7j�I���Y�}��u����Y�E��E������_   �]�;�t�uWS跙����;�uaVj�5<
����;�uL9=�t3V����Y���r����E;��P����    �E���3��uj�����Y�;�u�E;�t�    �������jh��蓳���]��u�u�����Y��  �u��uS襚��Y�  �=�#��  3��}�����  j�V���Y�}�S�����Y�E�;���   ;5�#wIVSP��������t�]��5V�k���Y�E�;�t'�C�H;�r��PS�u��-���S�u����E�SP������9}�uH;�u3�F�u������uVW�5<
���E�;�t �C�H;�r��PS�u��ٔ��S�u��I������E������.   �}� u1��uF������uVSj �5<
�������u�]j����YË}����   9=�t,V�����Y�����������9}�ul����P�U���Y��_����   �~���9}�th�    �q��uFVSj �5<
�������uV9�t4V����Y��t���v�V����Y�2����    3�����������|�����u��������P������Y����U����u�M��Ѵ���E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap���jj �t$j �������SVW�T$�D$�L$URPQQhXAd�5    ���3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�r/  �   �C�/  �d�    ��_^[ËL$�A   �   t3�D$�H3�赑��U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j��.  3�3�3�3�3���U��SVWj j h�AQ�k  _^[]�U�l$RQ�t$������]� U��QV�uV�9  �E�F��Yu�'���� 	   �N ����-  �@t����� "   ��S3ۨt��^��   �N�����F�F����f��F�^�]�u,�u7  �� ;�t�i7  ��@;�u�u��6  ��YuV�6  Yf�FW��   �F�>�H��N+�I;��N~WP�u�5  ���E��M�� �F����y�M���t���t������������#��0��@ tjSSQ�.  #����t%�F�M��3�GW�EP�u�35  ���E�9}�t	�N �����E%�   _[^���A@t�y t$�Ix��������QP�z���YY���u	���U��V����M�E�M�����>�t�} �^]��G@SV����t4� u.�D$�-��L$������C�>�u�\����8*u�ϰ?�i����|$ �^[�U��$�����x  ���3ŉ��  ��   S��  V3�W��  ��  �M��EЉ}ԉu��u�u��u��uĉu��u��ϰ��9u�u-�����VVVV�    V�@������}� t�E��`p������  �E��@@��   P��6  ���Yt6�u���6  ���Yt(�u���6  �u����4��#��6  ����YY3���0��@$�u����u��6  ���Yt6�u��6  ���Yt(�u��6  �u����4��#�o6  ����YY3���0��@$��"���;������3Ʉ҉ủu؉u��U���  C�}� �]���  ��, <Xw�������3��3�3����(�j��Y;��E��z  �$��M�M���u��u��u��uĉu�u��X  �� t>��t-��tHHt���9  �M��0  �M��'  �M��  �M�   �  �M��	  ��*u ���}ԋ�;��}���  �M��]���  �E�k�
�ʍDЉE���  �u���  ��*u���}ԋ�;��}���  �M���  �E�k�
�ʍDЉE��  ��ItF��ht8��lt��w�x  �M�   �l  �;luC�M�   �]��W  �M��N  �M� �E  �<6u�{4uCC�M� �  �]��(  <3u�{2uCC�e�����]��  <d�  <i��  <o��  <u��  <x��  <X��  �u��E�P��P�u���5  Y���E�Yt�MЍu�������C���]���  �MЍu�������  ��d�r  ��  ��S��   tZ��AtHHt@HHtHH�N  �� �E�   �U�M�@9u��]�   �]܉E���  �E�   �	  f�E�0uu�M�   �lf�E�0u�M�   �M����u������f�E��}ԋ��}���  ;�u�,��E܋E��E�   �  ��X�9  HHt]+��d���HH��  ��f�E��}�t'�G�Ph   �E�P�E�P�4  ����t�E�   ��G��E��E�   �E�E��P  ���;Ɖ}�t.�H;�t'f�E� � �M�t�+����E�   �  �u��  �(��E�P�H���Y��  ��p��  �t  ��e��  ��g�������itY��nt��o��  �E��E�   tI�M�   �@�7���}��d2  ����  �E� t	f�E�f���Ẻ�E�   �  �M�@�E�
   �M�f���C  ��W���k  u��guG�E�   �>9E�~�E��}�   ~-�u���]  V�8������U�Y�E�t
�E܉u�����E�   3�����E��G��E��E�P�u����u��}�P�u��E�SP�5�覗��Y�Ћ}����   t9u�u�E�PS�5$�耗��Y��YY�}�gu;�u�E�PS�5 ��a���Y��YY�;-u�M�   C�]�S�r����E�   �M��!��s�p���HH��������Y  �E�'   �E��E�   ������E�Q�E�0�E��E�   ����f�� ��������� t��@�}�t�G���G�����@�G�t��3҉}���@t;�|;�s�؃� �ځM�   f�E� ��ڋ�u3ۃ}� }	�E�   ��e���   9E�~�E����u!Eč��  �E��M������t$�EؙRPSW�J  ��0��9�]�����~M��N�̍��  +�Ff�E� �E؉u�tL��t�΀90tA�M܋M��0@�2If90t@@;�u�+E����;�u�(��E܋E��I�8 t@;�u�+E܉E؃}� ��   �E�@t%f� t�E�-��t�E�+��t�E� �E�   �]�+]�+]��E�u�uЍE�Sj �;������uċ}ЍE̍M��K����E�Yt�E�uWSj0�E��������}� �E�tQ��~M�u܉E���M�Pj���  P�E�FPF�}0  ����u9E�t�u��E̍��  ������}� Yu���M����M�P�E������Y�}� |�E�tWSj �E��������}� t�u������e� Y�]�����E�t$�M��}Ԋ��)����
����    3�PPPPP�$����}� t�E��`p��E̋��  _^3�[襅�����  ��^G�E�E/FiFqF�F�GU��W�}3�������ك��E���8t3�����_��U����u�M��X����E����   ~�E�Pj�u�/  ������   �M�H���}� t�M��ap��Ã=H u�D$����A���j �t$����YY�U���SV�u�M��ަ���]�   ;�sT�M胹�   ~�E�PjS�!/  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P�|.  ��YYt�Ej�E��]��E� Y��V���� *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�   ��$���o�����u�E���M�3��e���}� t�M��ap�^[�Ã=H u�D$�H���w�� �j �t$�����YY�U���(���3ŉE�SV�uW�u�}�M�菥���E�P3�SSSSW�E�P�E�P�9  �E�E�VP�.  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�������U���(���3ŉE�SV�uW�u�}�M������E�P3�SSSSW�E�P�E�P�r8  �E�E�VP�#3  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�P������U��WV�u�M�}�����;�v;���  ��   r�=�# tWV����;�^_u^_]鏴����   u������r*��$�TR��Ǻ   ��r����$�hQ�$�dR��$��Q�xQ�Q�Q#ъ��F�G�F���G������r���$�TR�I #ъ��F���G������r���$�TR�#ъ���������r���$�TR�I KR8R0R(R RRRR�D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�TR��dRlRxR�R�E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��S�����$��S�I �Ǻ   ��r��+��$��R�$��S�S(SPS�F#шG��������r�����$��S�I �F#шG�F���G������r�����$��S��F#шG�F�G�F���G�������V�������$��S�I �S�S�S�S�S�S�S�S�D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$��S�� TTT,T�E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_��U��MSV�u3�;�W�yu����j^�0SSSSS�c��������   9]v݋U;ӈ~���3�@9Ew�ɿ��j"Y�����;��0�F~�:�t��G�j0Y�@J;��M;ӈ|�?5|�� 0H�89t�� �>1u�A��~W�q���@PWV�������3�_^[]�U��Q�U�BS��VW��% �  ��  #ωE�B��پ   �%�� �ۉu�t;�t�� <  �(��  �$3�;�u;�u�Ef�M�X��L��<  �]����������M��E���ΉH�u��P������Ɂ���  �։P�t�M�_^f�H[��U���0���3ŉE��ES�]V�E�W�EP�E�P����YY�E�Pj j���u�����f��9  �uЉC�E։�EԉC�E�P�uV�������$��t3�PPPPP�������M�_�s^��3�[��|���������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j貆��Y�U��E�M%����#�������Vt1W�}3�;�tVV�B  YY��ռ��j_VVVVV�8�7�������_��u��P�ut	��A  ����A  YY3�^]Ã%�# �jh�������e� f(��E�   �#�E� � =  �t
=  �t3��3�@Ëe�e� �E������E������U���3�S�E��E�E�S�X��5    P��Z+�tQ�3���E�]�U�M�   ��U��E�[�E�   t�^�����t3�@�3�[��������#3��U��� SVW�I���3�9��E��]��]�]���   h�������;��y  �5�h��W��;��c  P萈���$��W����P�{����$��W����P�f������E�P虅����YYtSSSSS�������}�u,h��W��P�1���;�Y��th��W��P����Y�����M�;�ty9�tqP�p����5����c���;�YY��tV;�tR��;�t�M�Qj�M�QjP�ׅ�t�E�u3�E�P�0�����YtSSSSS�������}�r	�M    �D�M   �;��;E�t1P�����;�Yt&��;ÉE�t��;E�tP�ׇ��;�Yt�u��ЉE��5�过��;�Yt�u�u�u�u����3�_^[�ËD$S3�;�VWt�|$;�w����j^�0SSSSS�d��������=�t$;�u��ً�8tBOu�;�t��
BF:�tOu�;�u�躹��j"Y����3�_^[�U��SV�u3�9]Wu;�u9]u3�_^[]�;�t�};�w�{���j^�0SSSSS�����������9]u��ʋU;�u��у}���u�
�@B:�tOu���
�@B:�tOt�Mu�9]u�;�u��}�u�EjP�\�X�x��������j"Y���낋L$V3�;�|��~��u��^á���^��ʸ��VVVVV�    �+��������^ËD$��t���8��  uP�U}��Y�3��U��E�MSVW3��x�E3ۉx�EC���xt�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�@  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�  �EPSj �u���M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]�U��j �u�u�u�u�u�u�
�����]�U����ESV3ۋ���C��u�t�]tS�?  Y����  �t�Etj�%  Y����w  ����   �E��   j�  �EY�   #�tT=   t7=   t;�ub��M����@ ��{L�H��M�����{,�@ �2��M�����z�@ ���M�����z�0 ��0 ��������   ���   �E��   3��t����W�}�����D��   ��E�PQQ�$�P  �M��]��� �����������}�E�������T���]�����Au���3��E�����f�E�����;�}"+��]�t��u���m��]�t�M�   ��m�Hu���t�E����]��E������_tj�  Y�e���u��Et�E tj �  Y���3���^��[�ËD$��t~��裳��� "   �藳��� !   ÊD$� tj��t3�@ètj��tjX�������U��� 3���H�;Mtd@��|�3����E�t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E��  �E�P�h�������uV�:���Y�E�^�Ë�L��h��  �u(�y  �u�����E ����U��=@� u(�u�E���\$���\$�E�$�uj�3�����$]�茲��h��  �u� !   �  �EYY]�U������   ���3ĉD$|�u �EP�u��������u%�d$@�P�EP�EP�u�E �uP�D$P�������u�������=@� u+��t'�u �E���\$���\$�E�$�uP������$�P�#����$��  �u �p  �EYY�L$|3��p����]�QQ�D$���$�$YY�U��QQ�E�E�M�]��  ��������f�E��E���U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]ËM��  #�f;�uj��f���u�E�� u9Utj��3�]�U�����U����Dz3��   3�f�E�uc�E�� u9MtU�]��������Au3�@�3���e�E   �t�M�eJ�Et�f�e��;�tf�M ��EQQQ�$��������%Q���EQQ�$������U�����  �����  �E�]�Q��<$�$Y�Q�<$���$Y�U��Q��}��E�M#M��#E�����E�m�E���QQ�L$��t�-X �\$���t����-X �$������t
�-d �$���t	�������؛�� t���$�YY�jh���[���3�9�#tV�E@tH9p t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%p  �e��U�E�������e��U�;����U������   ���3ĉ�$�   �E�SV�u�HW�L$t+Ht$HtHtHtHHtHutj��   �hj�
j�j�j[Q�~WS�l�������uG�E��t��t��t�d$P���L$P�F����\$@���L$PW�NQPS�D$P�D$$P� �����h��  �t$�M����>YYt�=@� uV�������Yu�6�����Y��$�   _^[3��Bm����]��V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ����������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� j
j �t$�&8  ���V�t$����  �v�2r���v�*r���v�"r���v�r���v�r���v�
r���6�r���v ��q���v$��q���v(��q���v,��q���v0��q���v4��q���v��q���v8��q���v<�q����@�v@�q���vD�q���vH�q���vL�q���vP�q���vT�q���vX�q���v\�xq���v`�pq���vd�hq���vh�`q���vl�Xq���vp�Pq���vt�Hq���vx�@q���v|�8q����@���   �*q�����   �q�����   �q�����   �	q�����   ��p�����   ��p�����   ��p�����   ��p�����   ��p�����   ��p�����   �p����,^�V�t$��t5�;HtP�p��Y�F;LtP�p��Y�v;5PtV�zp��Y^�V�t$��t~�F;TtP�]p��Y�F;XtP�Kp��Y�F;\tP�9p��Y�F;`tP�'p��Y�F;dtP�p��Y�F ;htP�p��Y�v$;5ltV��o��Y^���U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^��U��QQ���3ŉE���SV3�;�W��u:�E�P3�FVh��V����t�5��4����xu
jX���������   ;���   ����   9]�]�u��@�E�5ذ3�9] SS�u���u��   P�u�֋�;���   ~<�����w4�D?=   w�`2  ��;�t� ��  �P�n��;�Yt	� ��  ���؅�ti�?Pj S�m����WS�u�uj�u�օ�t�uPS�u���E�S�����E�Y�u3�9]u��@�E9]u��@�E�u�U4  ���Yu3��G;EtSS�MQ�uP�u�{4  ����;�t܉u�u�u�u�u�u��;��tV�n��Y�Ǎe�_^[�M�3��h����U����u�M������u$�M��u �u�u�u�u�u�������}� t�M��ap�����U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^��U������3ŉE�SV3�9�W��u8SS3�GWh��h   S����t�=������xu
��   9]~"�M�EI8t@;�u�����E+�H;E}@�E������  ;���  ����  9] �]�u��@�E �5ذ3�9]$SS�u���u��   P�u �֋�;���  ~Cj�3�X����r7�D?=   w��/  ��;�t� ��  �P�k��;�Yt	� ��  ���E���]�9]��=  W�u��u�uj�u �օ���   �5�SSW�u��u�u�֋�;ˉM���   f�E t)9]��   ;M��   �u�uW�u��u�u���   ;�~Ej�3�X���r9�D	=   w�:/  ��;�tj���  ���P��j��;�Yt	� ��  �����3�;�tA�u�VW�u��u�u����t"9]SSuSS��u�u�u�VS�u �l��E�V�����Y�u�������E�Y�Y  9]�]�]�u��@�E9] u��@�E �u�1  ���Y�E�u3��!  ;E ��   SS�MQ�uP�u �-1  ��;ÉE�tԋ5�SS�uP�u�u��;ÉE�u3��   ~=���w8��=   w�$.  ��;�t����  ���P��i��;�Yt	� ��  �����3�;�t��u�SW��h�����u�W�u�u��u�u��;ÉE�u3��%�u�E��uPW�u �u��|0  ���u������#u�W����Y��u�u�u�u�u�u����9]�t	�u���i��Y�E�;�t9EtP��i��Y�ƍe�_^[�M�3���c����U����u�M������u(�M��u$�u �u�u�u�u�u�-����� �}� t�M��ap������U��SVWUj j h�o�u�>  ]_^[��]ËL$�A   �   t2�D$�H�3��Uc��U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h�od�5    ���3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y�ou�Q�R9Qu�   �SQ���SQ���L$�K�C�kUQPXY]Y[� ���U��QQ�EV�u�E��EWV�E��0  ���;�Yu�h���� 	   �ǋ��J�u�M�Q�u�P���;ǉE�u����t	P�Z���Y�ϋ������#�����D0� ��E��U�_^��jh�芀������u܉u��E���u������  ����� 	   �Ƌ���   3�;�|;�#r!�բ���8転��� 	   WWWWW�������ȋ������#��������L1��u&蔢���8�z���� 	   WWWWW�ۻ����������[P�0  Y�}���D0t�u�u�u�u�������E܉U���,���� 	   �4����8�M���M���E������   �E܋U�������u�B0  Y�U��$������  ���3ŉ�  ��   V3�9�$  �E��u��u�u3���  ;�u'�á���0詡��VVVVV�    �
���������  SW��  �����4��#�����ǊX$������u��]�t��u3��$  ����u&�Z���3��0�>���VVVVV�    蟺�����0  �@ tjj j ��  �~�������  �N  ��Y�9  ��D��,  �p���@l3�9H�E���P��4�M�������  3�9M�t����  ����]��E�3�9�$  �E��G  �E��E����=  ��u�3���
���E��ǃx8 t�P4��  ��	  �`8 j��  P�E��P�	  ��Yt4�M�+��$  3�@;��V  j�E�SP�a0  �������  C�E��jS�E�P�C0  �������  3�PPj��  Qj�M�QP�u�C�E��l������v  j �E�PV��  P�E�� �4������I  �E��M��9u��E��>  �}� ��   j �E�Pj��  P�E�� ƅ  �4�������  �}���  �E��E��a<t<u�33�f��
��CC�E��u��M�<t<u9�u��-  f;E�Y��  �E��}� tjXP�E��g-  f;E�Y��  �E��E���$  9E��H����  ���E��T4��D8�k  3ɋ��@��+  �ۋE��M���   9�$  �E��t  ��u��M��e� +M��E�;�$  s'�U��E��A��
u
�E�� @�E��@�E��}�   rы؍E�+�j �E�PS�E�P��4�������  �E�E�;���  �E�+E�;�$  r��  ���E���   9�$  ��  ��u��M��e� +M��E�;�$  s3�U��E��AAf��
u�E�f�  @@�E��E�f�@@�}��  rŋ؍E�+�j �E�PS�E�P��4������$  �E�E�;��  �E�+E�;�$  �p����  9�$  �2  �M��e� +M�j���  ^;�$  s,�U��u��f��
u
f�  �u�u�f�Ɓ}�R  r�3�VVh�  ��  Q���  +��+���P��PVh��  �l���;�tyj �E�P��+�P��5  P�E�� �4�����t	u�;���	���E�;�G�E�+E�;�$  �E��6����0j �M�Q��$  �u��0�����t�E��e� �E��	���E��}� u]�}� t'j^9u�u�;���� 	   �C����0�6�u��J���Y�+�u���D@t�E��8u3�������    �����  �����E�+E�_[��  3�^�Z����  ��jh(��Oy���E���u�͛���  貛��� 	   ����   3�;�|;�#r!褛���8芛��� 	   WWWWW�������ɋ������#��������L1��t�P��(  Y�}���D0t�u�u�u�?������E���'���� 	   �/����8�M���E������	   �E���x����u�D)  Y���h   �m����Y�L$�At�I�A   ��I�A�A�A   �A�a �ËD$���u襚��� 	   3��V3�;�|;�#r舚��VVVVV� 	   ������3�^Ëȃ������#���D��@^ø�á�#��Vj^u�   �;�}�ƣ�#jP�1m����YY�xujV�5�#�m����YY�xujX^�3ҹ���x��� ���� |�j�^3ҹ�W�������#����������t;�t��u�1�� B��|�_3�^��,  �=	 t��)  �5x�<^��Y�V�t$��;�r"�� w��+�����Q�����N �  Y^Ã� V���^ËD$��}��P�ō���D$�H �  YËD$�� P���ËD$��;�r= w�`���+�����P訌��YÃ� P���ËL$���D$}�`�����Q�~���YÃ� P���ËD$V3�;�u褘��VVVVV�    ���������^Ë@^á����3�9������U���SV�u3�;�W�}u;�v�E;�t�3���E;�t�������v�4���j^SSSSS�0薱�������R�u�M���x���E�9X��   f�Ef=� v6;�t;�vWSV�[��������� *   �ڗ��8]�� t�M��ap�_^[��;�t.;�w(躗��j"^SSSSS�0������8]�t��E��`p��u�����E;�t�    8]��0����E��`p��$����MQSWVj�MQS�]�p�l�;�t9]�b����M;�t�������z�H���;��k���;��c���WSV�JZ�����S���j �t$�t$�t$�t$�������U����u�M���w���E�M����   �A% �  �}� t�M��ap���j �t$����YY�U���S�u�M��w���]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�u�����YYt�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP������� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[��U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  �������W�M�E�u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5(N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r;�ur��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�$��+(;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5(N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��,A����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ; �,��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}� �4�3�@�   �4�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+,��M���Ɂ�   �ً0]���@u�M�U�Y��
�� u�M�_[��U���,�E�H
S�ف� �  �M�H�M��H� ���  ���?  �������W�M�E�u'3�3�9\��u@��|�3��  3��}૫j�X�  �e V�u��}ԥ���5@N�N���������с�  ��]��E�yJ���B�|��j3�Y+�@���M����   �E������҅T����|�� u@��|��n�ƙjY#������  �yN���F�e� +�3�B��L���1�u�19ur"9U���t+�e� �L����r;�ur��s�E�   H�U��M�yщM�M������!�E�@��}jY�|��+�3��} tC�<��+@;�}3��}૫��  ;��  +E��uԋȍ}ख़��¥������  ��yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�5@N�N���������с�  ��E�yJ���BjY+�3�B��\���M����   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e 3�+�B��L���1�<;�r;�s�E   �9�M���t�L����r3�;�r��s3�G�1��HyދM������!�E�@��}jY�|��+�3��DA����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�j3�X�Z  ;8�D��   3��}૫��M�   �����������  �yJ���B�e� �e ��������E�    )U��׋]�\���3��#ωM�����M�u�3�u����E�}�u�|Ӌ�j���M�Z+�;�|�1�t����d�� J����}�8�L�3�@�   �L�e����؋���������  �yJ���B�e� �e ��������E�    )U��֋M�|����#ΉM�����M}�|���}��M����E�}�}�|Ћ�j���M�Z+�;�|�1�t����d�� J����}�3�^jY+D��M���Ɂ�   �ًH]���@u�M�U�Y��
�� u�M�_[��U���|���3ŉE��ES3�V3��E��EF3�9]$W�E��}��]��u��]��]��]��]��]��]��]�u�+���SSSSS�    茤����3��  �U�U��< t<	t<
t<uB��0�B���/  �$�w��Ȁ�1��wjYJ�݋M$�	���   �	:ujY������+tHHt����  ���jY�E� �  뢃e� jY뙊Ȁ�1���u�v��M$�	���   �	:uj�<+t(<-t$:�t�<C�<  <E~<c�0  <e�(  j�Jj�y����Ȁ�1���R����M$�	���   �	:�T���:��f����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�]���<+t�<-t��`����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*�<	�u��n���j�����J��M��Ȁ�1��wj	��������+t HHt���;���j�����M��jY�@���j�o����u���B:�t�,1<v�J�(�Ȁ�1��v�:�뽃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�[����B:�}��O����M��E�O�? t�E�P�u��E�P��  �E�3Ƀ�9M�}��E�9M�uE9M�u+E=P  ��  =������  ���`;��E���  }�ؾh�E���`9Muf�M�9M���  �E��}���T�����u��q  k�Ƌ�f�; ��]�r��}�����M��u��]��]��S
�M�3��E��EԉE؉E܋¿�  3�#�#�% �  f����<
����  f�����  f������  f���?w3��EȉE���  f��uG�E����u�}� u�}� u	f!M���  3�f;�u!G�C���u9Ku9u�M̉MȉM��  !M��u��E�   �M��U�Ʌ҉U�~U�Lă��M��]��M��U���	�e� �ʋV��
;�r;�s�E�   �}� �^�tf��E��m��M��}� ��]�FF�E��M��}� ����  f��~;�E�   �u-�u؋M��e�������M����ʁ���  f���u؉M��f��M����  f��}B��������E�t�E��M܋]؋U��m�����ًM������N�]؉M�u�9u�tf�M�f�}� �w�Mԁ��� �� � u3�}��u*�e� �}��u�e� f�}���u	f�E� �G�f�E���E���E�f����u�sf�M�f�MċM؉MƋM���M�f�}��f����e� %   � ���e� �Ẽ}� �m����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W�M�_^3�[�C�����Ӊ)�\���ي�H�3�����V�U���t���3ŉE�S�]VW�u�}�f��U��ʸ �  #ȁ��  f�ɉ]��E���E���E���E���E���E���E���E���E���E���E���E�?�E�   �M�t�C-��C f�ҋu�}�u.��u*��u&f!;f;�����$ �C�C�C0�C 3�@��  f�����   �   �;�f� u��t��   @uh���Qf��t��   �u��u;h���;�u0��u,h���CjP�;�����3���tVVVVV�������C�*h���CjP������3���tVVVVV�ܛ�����C3��  �ʋ�i�M  �������Ck�M���������ىM�3���ۃ�`;�f�U�u�}�f�E��M���  }�h�ۃ�`�M�;���  �E�T�˃������y  k�M�f�9 ��M�r��}ĥ��Eĥ�MƉE����y
�U�3��Ͼ�  3�#�#��E��E��E�E��� �  f;֍���  f;���  f=����  f=�?w3��E�E�E���  3�f;�u@�E����u9u�u9u�u	f�u���  f;�u$�U�@�B���u9ru92u�u�u�u��  �}�u��}��E�   �U��u�҅��u�~X�T��U��U����U��U��u��6����փe� �4;�r;�s�E�   �}� �}��w�tf��E��m��M��}� �GG�E��M��}� �}���  f��~;�E�   �u-�U��}�u��e������U�������  f���}�U��f��R��  f��}H�����҉U���E�t�E��U��}�u��m�������U�������M��}�U�uσ}� tf�M�f�}� �w�U����� �� � u3�}��u*�e� �}��u�e� f�}���u	f�E� �@�f�E���E���E�f=�sf�U�f�U��U�U�U���U�f�E��f��Ƀe� ��   ��� ���e� �M���k���3��M���f���?��  �H  �u��E��ы�3�#�#�� �  f;Ӎ<�E��E��E�E�����  f;���  f������  f���?w�E���  f;�uG�E����u9E�u9E�u	f�E���  f;�uG�E����u
9E�u9E�t��e� �E��E�   �U��u�҅��u�~R�u؍T��u��U��U��u��6��e� �֋p��;�r;�s�E�   �}� �X�tf� �E��m��M��}� �@@�E��M��}� ����  3�f;�~<�E�   �u.�U��]�u��e����ڋU����ց���  f;��]�U��f;�M����  f;�}B��������E�t�E��U��]�u��m�����ڋU������H�]�U�u�9E�tf�M�f�}� �w�U����� �� � u1�}��u(�}���E�uf�}����E�u	f�E� �G�f�E���E���E�f���rf�ىE�E�Ɂ�   ��� ���M�3��6f�E�f�E��E�E�E���E�f�}���f��Ɂ�   ��� ���M�E�E��E�U��M�f�
t2��M9E'f�" f�}� ��B����$ �B�B0�B ����jY9M~�M�u���j���?  f�E�[�E��}�M��e������E�����K�}�E�uڅ�}2�ށ��   ~(�E�}�M��m�������E������N���}�E�؋E@���Z�]��E���   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B�ҋ�tA�Eȍ0;։U�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K���K�K<5}�M��D�;9u	�0K;]�s�;]��E�sCf� �*؀��ˈX�D �E��M�_^3�[��:���À;0uK;�s�;ًE�s�f�  f�}� ��@���ʀ��� �P�0�@ �����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u�����   ^t   �3���t��   ��SVW�   t���t   ��t   ��t   ��   �   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#с�   ^[t��   t
;�u �  Ã�@�@�  Ã�SUVW��|$�\$3���tjZ��t����t����t���� t����t��   �ˋ��   #ǽ   �   t =   t=   t;�u��
����   #�t;�u��   ���   f�� t��   �t$(�L$$����#�#��;D$��   ���������D$�l$��|$�\$3���tjZ��t����t����t���� t����t��   �ˋ�#�t$=   t=   t;�u����   ���   #�t��   u��   ���   f�� t��   �T$�=�# ��  �����\$�D$3���yj^f� t��f� t��f� t��f� t��f� t��   �Ƚ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #Ã�@t-�  t��@u��   ���   ���   ��#|$$��#��;�u���   �"���P�D$,����Y�\$(�D$(3҄�yjZ�   ��t��f� t��f� t��f� t���   ��t��   ��#�t"��    t�� @  t;�u��   ����#Ã�@t-�  t��@u��   ���   ���   �L$��3���� t   �_^][�����Q�L$+ȃ����Y��  Q�L$+ȃ����Y��  U���VW�u�M��gX���E�u3�;�t�0;�u,�jw��WWWWW�    �ː�����}� t�E�`p�3���  9}t�}|Ƀ}$ËM�S��}��~���   ~�E�P��jP�[����M������   ���B����t�G�ǀ�-u�M���+u�G�E���I  ���@  ��$�7  ��u*��0t	�E
   �4�<xt<Xt	�E   �!�E   �
��u��0u�<xt<XuG�G���   ���3��u���N��t�˃�0�f��t1�ˀ�a����w�� ���;Ms�M9E�r'u;�v!�M�} u#�EO�u �} t�}�e� �\�]��]ى]��G댨����u�u>��t	�}�   �w	��u,9u�v'��u���E� "   t�M����E$�����ƉE��E��t�8�Et�]��}� t�E�`p��E���E��t�0�}� t�E�`p�3�[_^��U��3�9HP�u�u�uuh ��P������]�U������3ŉE�j�E�Ph  �u�E� �ܰ��u����
�E�P�j���Y�M�3���3����U���4���3ŉE��E�M�E؋ES�EЋ V�E܋EW3�;E�M̉}��}��_  �5İ�M�QP�օ��ذt^�}�uX�E�P�u�օ�tK�}�uE�u܃���E�   u�u��t�����YF;�~[�����wS�D6=   w/������;�t8� ��  �-WW�u��u�j�u�Ӌ�;�u�3���   P�8��;�Yt	� ��  ���E���}�9}�t؍6PW�u��,7����V�u��u��u�j�u�Ӆ�t�]�;�tWW�uSV�u�W�u�l���t`�]��[9}ԋl�uWWWWV�u�W�u�Ӌ�;�t<Vj�F��;�YY�E�t+WWVPV�u�W�u��;�u�u��28��Y�}���}��t�MЉ�u�諺��Y�E��e�_^[�M�3��2���ËL$S3�;�VW|[;�#sS������<��#�������@t5�8�t0�=�u+�tItIuSj��Sj��Sj�� ����3����r��� 	   ��r������_^[ËD$���u��r���  �r��� 	   ����V3�;�|";�#s�ȃ������#����@u$�r���0�qr��VVVVV� 	   �ҋ�������^Ë ^�jhH���O���}����������4��#�E�   3�9^u6j
�f��Y�]�9^uh�  �FP�I���YY��u�]��F�E������0   9]�t�����������#�D8P����E��O���3ۋ}j
�te��YËD$�ȃ������#���DP����U������3ŉE�V3�95 tN�=D�u�K  �D���uf���pV�M�Qj�MQP����ug�= u�����xuЉ5 VVj�E�Pj�EPV��P�l��D���t�V�U�RP�E�PQ����t�f�E�M�3�^�/�����    ��U���SV�u3�;�t9]t8u�E;�tf�3�^[���u�M��Q���E�9Xu�E;�tf�f�8]�t�E��`p�3�@�ʍE�P�P�q�����YYt}�E����   ��~%9M| 3�9]��R�uQVj	�p�ذ���E�u�M;��   r 8^t8]����   �e����M��ap��Y�����o��� *   8]�t�E��`p�����:���3�9]��P�u�E�jVj	�p�ذ���:����j �t$�t$�t$��������jhh��#M��3ۉ]�j�$d��Y�]�j_�}�;=�#}W�����x�9tD� �@�tP��  Y���t�E��|(�x��� P�X��x�4��3��Y�x�G��E������	   �E���L���j��b��Y�SV�t$�F�Ȁ�3ۀ�u?f�t9�FW�>+���~,WPV�%���YP�������;�u�F��y����F��N ���_�F�f �^��[�V�t$��u	V�3   Y^�V������Yt���^�f�F @tV�����P�  YY���^�3�^�jh����K��3��}�}�j��b��Y�}�3��u�;5�#��   �x��98t^� �@�tVPV�����YY3�B�U��x���H���t/9UuP�P���Y���t�E��9}u��tP�5���Y���u	E܉}��   F�3��u�x�4�V�����YY��E������   �}�E�t�E��aK���j�Ia��Y�j����Y�U������3ŉE��ESV3�9uW�E�N@  �0�p�p�F  ��X���}𥥥�����<�ыH�����Ή}���e� �������ˋ]���׍<;��0�P�Hr;�s�E�   3�9]�8t�r;�r��s3�C�ۉptA�H�H�U�3�;�r;�s3�F���Xt�@�M�H�e� �?�����<��P������Uމ�x�X��4;�U�r;�s�E�   �}� �0t�O3�;�r��s3�B�҉HtC�X�M�E�} �����3��&�H�����P�����������E���  �H�9ptջ �  �Xu0�0�x�E���  ������0�4?�H�����ʅˉp�Ht�f�M�f�H
�M�_^3�[�*���������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � �������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_��3�PPjPjh   @h����DáD���V�5�t���tP�֡@���t���tP��^�SV�t$W3����;�u�j��WWWWW�    ��������B�F�t7V����V����  V�����P�  ����}�����F;�t
P�*/��Y�~�~��_^[�jh����G���M��3��u3�;���;�u�<j���    WWWWW蝃���������F@t�~�E���G���V����Y�}�V�/���Y�E��E������   �ՋuV�����Y�jh���aG���E���u��i��� 	   ����   3�;�|;�#r�i��� 	   SSSSS�������Ћ����<��#��������L��t�P����Y�]���Dt1�u����YP����u���E���]�9]�t�Ji���M��-i��� 	   �M���E������	   �E���F����u�Q���Y�V�t$WV�2������YtP����#u	���   u��u�@Dtj����j�������;�YYtV�����YP����u
�����3�V�S����������#������Y�D0 tW�h��Y����3�_^�jh����E���E���u�gh���  �Lh��� 	   ����   3�;�|;�#r!�>h���8�$h��� 	   WWWWW腁�����ɋ������#��������L1��t�P����Y�}���D0t�u�����Y�E����g��� 	   �M���E������	   �E��xE����u�����Y�V�t$�F��t�t�v�D,���f����3�Y��F�F^����̍B�[Í�$    �d$ 3��D$S�����T$��   t�
��:�tτ�tQ��   u��W����V؋
����~����3���������3�3ƃ��� �u% �t�% u��   �u�^_[3�ËB�:�t6��t�:�t'��t���:�t��t�:�t��t��^_�B�[ÍB�^_[ÍB�^_[ÍB�^_[��%԰������������h��.��Y����̃=p uK�h��t�`�Q<P�B�Ѓ��h    �t��tV���0f��V��������t    ^�                                                                                                                                                                                                                                                                                                                                                                                                                                                                           T� j� |� �� �� �� �� �� �� �� �� � � "� ,� D� T� l� t� �� �� �� �� �� �� �� � 0� F� `� n� |� �� �� �� �� �� �� � (� F� Z� f� ~� �� �� �� �� �� �� �� � �  � ,� B� T� f� x� �� �� �� �� �� �� �� �� � $� 2� @�         Э        ��'=zXz        `��z            bad allocation  ||----------------------------------------  ||  http://www.biomekk.com  ||  (c) 2009 Christopher Montesano  $�P" p  �l `! �l �l �l �l t�p! 0 � �� ��    �� �� ��     0�P" �! �l `! �l �l �l �l select_nth.tif  c:\program files\maxon\cinema 4d r12\plugins\selectloop\source\selectloop_cmd.h .00 .0  ||   - ERROR: Component Initialization Failed   ||   - Component Successfully Loaded    ||       v  select_loop.tif     c:\program files\maxon\cinema 4d r12\resource\_api\c4d_general.h    %s                 ����MbP?��g PL ���f     c:\program files\maxon\cinema 4d r12\resource\_api\c4d_baseobject.cpp   H�@l res          �f@-DT�!	@      �?\��� `� p� �� �� �� �� �� �x       Y@     @�@p��� `� p� �� �� �� �� �� �� ��P� 0� @� е � P� �� � ��  � � c:\program files\maxon\cinema 4d r12\resource\_api\c4d_gui.cpp  ���� `� p� �� �� �� �� �� � ��� `� p� �� �� �� �� �� �� �  � 0� @� P� `� p� `� �� �� �� �� Progress Thread 0%  ~   %       c:\program files\maxon\cinema 4d r12\resource\_api\c4d_resource.cpp #   M_EDITOR        c:\program files\maxon\cinema 4d r12\resource\_api\c4d_file.cpp �������������      �?c:\program files\maxon\cinema 4d r12\resource\_api\c4d_libs\lib_ngon.cpp        c:\program files\maxon\cinema 4d r12\resource\_api\c4d_basebitmap.cpp   c:\program files\maxon\cinema 4d r12\resource\_api\c4d_basetime.cpp      �Ngm��C   ����A  4&�k�  4&�kCh��z�z����    c:\program files\maxon\cinema 4d r12\resource\_api\c4d_pmain.cpp    ��P�    c:\program files\maxon\cinema 4d r12\resource\_api\c4d_gv\ge_mtools.cpp ����@�0���������    �n�n�              �?      �?3      3            �      0C       �       ��              CorExitProcess  mscoree.dll .mixcrt EncodePointer   KERNEL32.DLL    DecodePointer   FlsFree FlsSetValue FlsGetValue FlsAlloc    e+000      �~PA   ���GAIsProcessorFeaturePresent   KERNEL32    @
�
runtime error   
  TLOSS error
   SING error
    DOMAIN error
      R6034
An application has made an attempt to load the C runtime library incorrectly.
Please contact the application's support team for more information.
      R6033
- Attempt to use MSIL code from this assembly during native code initialization
This indicates a bug in your application. It is most likely the result of calling an MSIL-compiled (/clr) function from a native constructor or from DllMain.
  R6032
- not enough space for locale information
      R6031
- Attempt to initialize the CRT more than once.
This indicates a bug in your application.
  R6030
- CRT not initialized
  R6028
- unable to initialize heap
    R6027
- not enough space for lowio initialization
    R6026
- not enough space for stdio initialization
    R6025
- pure virtual function call
   R6024
- not enough space for _onexit/atexit table
    R6019
- unable to open console device
    R6018
- unexpected heap error
    R6017
- unexpected multithread lock error
    R6016
- not enough space for thread data
 
This application has requested the Runtime to terminate it in an unusual way.
Please contact the application's support team for more information.
   R6009
- not enough space for environment
 R6008
- not enough space for arguments
   R6002
- floating point support not loaded
    Microsoft Visual C++ Runtime Library    

  ... <program name unknown>  Runtime Error!

Program:              �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow       �?5�h!���>@�������             ��      �@      �                    �������             ��      �@      �         Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ()  ,   >=  >   <=  <   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>  =    delete  new    __unaligned __restrict  __ptr64 __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(        ��������������|�p�d�(�����|�\�@�\�T�P�L�H�D�@�<�8�,�(�$� ���������� ���������|�������������������������������������t�h�T�4����������t�P�0������������������x�\�<��������|�X�4������(�InitializeCriticalSectionAndSpinCount   kernel32.dll    	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx          GetProcessWindowStation GetUserObjectInformationA   GetLastActivePopup  GetActiveWindow MessageBoxA USER32.DLL  _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh                                                                                                                                                                                                                                                                                          ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun     1#QNAN  1#INF   1#IND   1#SNAN  SunMonTueWedThuFriSat   JanFebMarAprMayJunJulAugSepOctNovDec    CONOUT$ ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           �� �              ������    �       ����    @   �� �        ����    @   �           ���                8�8�           H�X�����    8�       ����    @   8�            X���           ��������    X�       ����    @   ��x�       ����    @   ��           ������    ��        ����    @   �           (���                ��D�           T�d�����    ��       ����    @   D�           ����    ��        ����    @   ��            ����           ����    ��        ����    @   ��            ��            �,���    �       ����    @   �             ��            ���            x���            D���           ����    D�        ����    @   ��            `���           ������    `�       ����    @   ��            x�,�           <�L�����    x�       ����    @   ,�            ��|�           ����    ��        ����    @   |�            ����           ����    ��        ����    @   ��            ��           �$�    �        ����    @   �            4�T�           d�p���    4�       ����    @   T�            X���           ����    X�        ����    @   ��            ����           �� �    ��        ����    @   ��    P� XA �o                     ����    ����    ����k�|�    ����    ����    ����    P�    ����    ����    ����    r�    ����    ����    ����    ��    ����    ����    ����    i�    ����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    $�����    0�����    ����    ����9�=�    ����    ����    ����    �    ����    ����    ����    �    ����    ����    �����/0    ����    ����    ����K0O0    ����    ����    ����    =2    ����    ����    ����)3@3    ����    ����    ����    b6    ����    ����    ����    9    ����    ����    ����    �<    ����    ����    ����    ">    ����    ����    ����    �?    ����    ����    �����WX    ����    ����    �����d�d    ����    ����    ����    ar    ����    ����    ����    _y    ����    ����    ����    ��    ����    ����    ����    O�    ����    ����    ����    ͦ        ������    ����    ����    p�    ����    ����    ����    R�    ����    ����    ����    ��4�         T�  �                     T� j� |� �� �� �� �� �� �� �� �� � � "� ,� D� T� l� t� �� �� �� �� �� �� �� � 0� F� `� n� |� �� �� �� �� �� �� � (� F� Z� f� ~� �� �� �� �� �� �� �� � �  � ,� B� T� f� x� �� �� �� �� �� �� �� �� � $� 2� @�     FGetCurrentThreadId  GetCommandLineA HeapFree  �GetVersionExA HeapAlloc �GetProcessHeap  qGetLastError  �GetProcAddress  GetModuleHandleA  � ExitProcess eTlsGetValue cTlsAlloc  fTlsSetValue dTlsFree ,InterlockedIncrement  (SetLastError  (InterlockedDecrement  VSleep $SetHandleCount  �GetStdHandle  fGetFileType �GetStartupInfoA � DeleteCriticalSection }GetModuleFileNameA  � FreeEnvironmentStringsA UGetEnvironmentStrings � FreeEnvironmentStringsW �WideCharToMultiByte WGetEnvironmentStringsW  HeapDestroy HeapCreate  �VirtualFree �QueryPerformanceCounter �GetTickCount  CGetCurrentProcessId �GetSystemTimeAsFileTime ^TerminateProcess  BGetCurrentProcess nUnhandledExceptionFilter  JSetUnhandledExceptionFilter 9IsDebuggerPresent �WriteFile QLeaveCriticalSection  � EnterCriticalSection  �VirtualAlloc  HeapReAlloc HeapSize  RLoadLibraryA  #InitializeCriticalSection GetCPInfo � GetACP  �GetOEMCP  ?IsValidCodePage �RtlUnwind uMultiByteToWideChar tGetLocaleInfoA  �RaiseException  �GetStringTypeA  �GetStringTypeW  DLCMapStringA  ELCMapStringW  SetFilePointer  "GetConsoleCP  3GetConsoleMode  7SetStdHandle  �WriteConsoleA 5GetConsoleOutputCP  �WriteConsoleW S CreateFileA 4 CloseHandle � FlushFileBuffers  KERNEL32.dll                    K?eL    ��          �� �� �� �� ��   selectloop.cdl c4d_main                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       `��    .?AVCommandData@@   �    .?AVBaseData@@  �    .?AVSelectNthCommand@@  �    .?AVSelectNthDialog@@   �    .?AVGeModalDialog@@ �    .?AVGeDialog@@  �    .?AVSelectLoopCommand@@ `�`�`��    .?AVGeSortAndSearch@@   �    .?AVNeighbor@@  �    .?AVDisjointNgonMesh@@  `�`�`�`�`��    .?AVGeUserArea@@    �    .?AVSubDialog@@ �    .?AViCustomGui@@    `�`�`�`�`�`�`�`�`�`�`�`��    .?AVC4DThread@@ `�`�`�`�`�`�`��    .?AVGeToolNode2D@@  �    .?AVGeToolDynArray@@    �    .?AVGeToolDynArraySort@@    �    .?AVGeToolList2D@@  `�`�`�`��    .?AVtype_info@@ u�  s�  N�@���D    sqrt            fmod         ���?��?�==g=��?�`�            ����������    �����
                                                                   �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �             x   
   OWOWOWOWOWOWOWOWOWOW          h�   <�	   �
   x�   L�   �   ��   ̼   ��   l�   4�   ��   Ի   ��   P�    �!    �"   ��x   l�y   \�z   L��   H��   8�                                                                                                                                                                                                                                                                                                                   	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                 ?             ���5�h!����?      �?             
      p?  �?   _       
          �?      �C      �;      �?      �?      ���d j o u z � � � � � � � � � � !!>!C!]!b!�!�!�!�!�!�!""&":"R"f"�"�"�"�"�"�"�"
#*#/#I#N#n#�#�#�#�#�#�#�#$&$>$R$r$w$�$�$�$�$�$  t�    C                                                                                              �            �            �            �            �                              H        p���x��  �    ��                                                                                                                                                                                                                                                                                                                                    abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                     ��  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��     ������            �&         ��   ��   ��   ��   d�   \�!   T�   ��   ��   ��   L�   D�   p�   l�    h�   ��   |�   <�   t�   4�   ,�   $�   �   �"   �#   �$   �%    �&   ��      �      ���������              �       �D        � 0                 p�r�����������������x�p�d�X�P�D�@�<�8�4�0�,�(�$� ����� �����0�����������������������x�	         � .   D���������H   .               �            �    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ���5      @   �  �   ����             �p     ����    PST                                                             PDT                                                             `�����        ����                        �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
            ����   ;   Z   x   �   �   �   �     0  N  m  ����   :   Y   w   �   �   �   �     /  M  l          ��������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             0040E0t0�0�0�0�0�0�0141I1[1l1~1�1�1�1�1�1�1�1�23X3s3�5\6�6�6�6�6�6�6�6	7E7W7�7�7�7�7�7�7�7848C8U8g8x8�8�8�8�8�899&9D9Y9k9}9�9�9�9�9�9�9�9�9:$:8:Q:c:x:�:�:�:�:�:;;&;8;J;d;v;�;�;�;�;�;�;�;	<4<F<X<_<|<�<�<�<�<�<:=M=y=�=�=O>a>�>�>�>�>�>??9?�?      �   ,0�0�0�1�2�2�2�2�2�23$3Q3d3�3�3�34$4T4�4�4�4545T5�5�5�5�56$6D6d6v6�6�6�6�6�67$7D7d7�7�7�78$8D8d8�8�8�8�8�8�8949T9t9�9�9�9:$:D:a:t:�:�:�:;;4;�;�;�;�;<4<T<t<�<�<�<�<=4=t=�=�=#>s>�>�>!?D?t?�?�?�? 0    0$0A0Q0d0�0�0�0�0191M1�1�1�1242T2t2�2�2�2�2$3B3V3f3�3�3�3�3444`4t4�4�4�4�45:5m5{5�5�5�5�5�56$6>6R6b6�6�6�6�67,7U7�7�7�7�7�7�7%8S8i8w8�8�8�899T9}9�9�9�9:4:_:�:�:�:�:;$;A;T;t;�;�;�;<$<D<d<�<�<�<�<=$=A=Q=d=�=�=�=�=�=>)>;>U>f>x>�>�>�>?$?T?�?�?�?�?   @  �   040a0�0�0�0141~1�1�12$2D2d2�2�2�23!3A3d3�3�3�3444d4�4�4�4�4515D5a5�5�5�5$6�6�6�6�6747d7�7�7�7818Q8q8�8�89$9D9t9�9�9�9$:d:�:�:;A;a;�;�;�;<$<2<7<T<}<�<�<*=T=t=�=�=>W>�>W?�?�?�?�? P  �   040]0�0�0�0$1A1d1�1�1�1�2�2�23$3T3�3�3�3�3444R4s4�4�4�4545Q5t5�5�5616T6�6�6�6�6!747T7�7�7818T8t8�8�8�89a9~9�9�9�9:2:[:l:�:�:�:�:;&;N;b;�;�;�;<%<[<s<�<�<�<�<�<�=�=>>W>_>�>�> `  �   �0�3�34-4f4v4�4�45�6�6�6�67 7Q7d7�7�7�7�7818T8t8�8�8�89$9A9d9�9�9�9T:�:�:;!;1;D;�;�;�;�;�;<$<L<�<�=�=�=�=�=�=�=�=>%>Y>?�?�? p  �   0<0d0�0�01%1�1�1	2%2�2�2	3,3H3l3�3�3�3�3M4e4�4<5a5�5�56$6D6d6q6�6�6�67$7�7�7�7�7<8h8�8�8�89W9%:*:5:Z:b:�:�:�:�:!;T;�;�;<D<k<�<�<
=6=K=t=�=�=+>k>�>�> ?d?�?�?�?�?   �  �   0'0V0m0�0�0�0121Q1p1�1�1�1202O2�2�2�2�23'3g3�3�3�3�3*4�4�4%5~5�56[6�6�6�6;7|7�7�7�7<8V8�8�89!9x9�9�9�94:�:;t;�;�;6<H<�<�<===�=�=->f>�>�>�>?/?F?t?�?�?�? �  t   0i01I1�1�132�2�2#3�3�3C4�4�4C5�56c6�6#7�7�7C8�8�8S9�9:�:�:);s;�; <:<`<�<�<�<$=N=�=�=>;>C>t>�>�>?Z?�?�? �  �   N0�0�01D1�1�1�12D2�2�2�213a3�3�3�3414�4�4�4�45"5�5�5�5�6V7�7�7�7�7�7�7�7�7�7�7�8 99999999 9�9�9�9:?:R:n:�:�:�:�:;4;d;�;�;�;<4<t<�<�<=1=|=�=$>D>d>�>�>�>?D?t?�?�?�?�?�?   �  �   0#070T0d0�0�0�0�0�0�01"1?1K1V1t1�1�1!2A2d2�2�2 3p3�3�3�3F4t4�4�45T5n56D6�6�6�6�6`7�7�7�7�7�8�8X9�9�9�9�9�9�9�9A:�:�:�:�:
;;D;d;�;(<�<	=4=d=�=�=�=->�>?!?T?t?�?�?�?�?   �  �   040d0�0�011)1H1Q1�1�1�1�23E3W3s3�3�3�3 4!4=4\4x4�4�4�45 5�5�5�5�5�516?6R6p6�6�6�6�6�67'7D7�7�7�78C8�8N9z9�9�9�9:D:r:�:�:;T;u;�;�;�;�;�;�;<+<K<x<�<�<�<�<�<�<�<=$=5=H=`=r=�=�? �  �   .0d0�01i1�1D2e2�2�2d3�3494�4	5�5�5�5	66,6<6Y6�6�6�6	7=7�7�7�7�7�78#8D8\8�8�8�8�8�8\:c:�:�:;';d;�;�;�;<<W<�<�<�<�<$=-=:=T=a=n=�=�=�=�=�=�=�=>'>B>X>t>�>�>�>�>�>�>	??-???H?f?�?�?�?�?�?�? �     00/0P0f0�0�0�0�0�0�011+1=1O1X1v1�1�1�1�1�122!2?2`2v2�2�2�2�2�2�23?3d3r33�3�3�3�3�3�34$464R4h4�4�4�4�4�4�45"545F5O5m5�5�5�5�5�56666L6w6�6�6�6R7Z7d7v7�7�7�7�7�7�7�7O8m8�8�8�8E9W9h9q9�9�9�9:4:H:Z:l:�:�:�:�:�;�;�;!<a<�<�<�<�<=$=T=f=�=�=�=�=$>D>a>�>�>�>�>?$?T?o?�?�?�?�? �  �   0$0T0�0�0�0�0141d1�1�1�12$2Q2t2�2�2�2343T3t3�3�3�3�3414D4d4�4�4�4.5N5c5�56a6�6�6X7z7�78:8]8�8�89~9�9�93:\:�:�:�:$;�;�;<�<�<�<c=�=�=.>N>c>�>L?w?�?�?   �   Q0w0�0�0Q1�132\2�2�2333�3�3�374�4�4l5�5�5�5�5�5$6D6[6�6�6�6�617Q7t7�7�7�7�7'8Q8�8�8�8�89+9J9�9�9�9�9:1:Q:t:;;;;?;a;�;�;�;�;<$<T<�<�<�<�<=!=1=U=�=�= >.>g>�>�>�>1?      �0�0�0+1�1�1�1�1�1�1�1�1�1�1�1�12222 243a3r3�3�3�3�3�3�34%434Q4b4�4�4�4�4�45,5@5P5t5�5�5�5�5�5�56,6@6O6_6p6�6�6�6�67$7D7d7�7�7�7�7�7848T8�8�8�8�8�8!949d9�9�9�9�9�9:1:A:Q:d:�:�:�:�:;$;D;d;�;�;�;�;�; <(<<<�<�<=!=E=�=�=�=�=>$>D>d>�>�>�>�>?!?1?D?q?�?�?�?�?�?�?     ,  0#010@0a0�0�0�0�0�011!141T1o1}1�1�1�1�1�1242T2t2�2�2�2�2'3@3Q3m3�3�3�3�3�3	444T4t4�4�4�4�455.5>5P5t5�5�5�5�5�5�56>6U6l6}6�6�6�6�6�67"767E7U7f7�7�7�788$8D8d8�8�8�8�89$9D9d9�9�9�9�9:$:D:d:�:�:�:�:;,;T;�;�;�;�;<$<D<d<�<�<�<�<=$=D=d=�=�=�=�=>$>D>d>�>�>�>�>�>?4?T?q?�?�?�?�?�?�?   0 �   060J0Z0�0�0�0�0�0�021G1�1�1�12$2t2�23T3t3�3�3�3�3444T4�4�4�4�4545a5�5�5�5616T6�6�6�6717Q7q7�7�7�7�7818Q8q8�8�8�8�8919Q9 @ $   �3A=a=�=�=>E>�>�>?R?�?�?�? P p   20e0�0�0%1b1�1�1�1"2U2�2�2%3u3�3�354u4�4%5�5h7�70:�:�:�:�:�:�;�;�;�;R<`<�<�<N=\=�=�=�=�=�>�>??�?�?�?�? ` �   �0�0�0�01$1T1�1�1�1�12$2T2�2�2�2�2343d3�3�3�3�344t4�4�4�4�4545T5�5�5�5�5q6�6�6�67$7�8
99@9�:1;D;t;�;�;�;<#<D<d<�<�<�<==$=Q=q=�=�=�=�=$>?<?�?�? p �   0�0�0�0�1�1�12a2k2�2373W3�3'4e4|4�4�4�45(5F5T5�5�5616T6q6�6�67e7q7{7�7�7�7�7�7�7,8Q8d8�8�8�8�89.989C9H9t9�9�9�9:A:a:�:�:�:;�;<B<u<�<�<%=u=�=�=>E>�>�>?_?�?�? � �   "0R0�0�01b1�1�1"2U2�2�2353e3�34E4�4�45#5P5d5t5�5�5%6e6�6�657u7�7898a8�8�8�8�8�89<9e9�9�9�9(:O:�:�:�:5;];�;�;�;"<V<x<�<U=r=�=�=�=�=>$>D>a>q>�>�>�>�>�>�>?4?T?t?�?�?�?�?   � �   0D0d0�0�0�0�01$1D1�1�1�1�1�12!2?2a22�2�2�2313T3t3�3�3�3�34$4A4T4t4�4�4q5�5�56K6�67U7�7�7&8u8�8�8(9�9�9:E:�:�:;X;�;�;"<U<�<�<�<E=�=�=�=�=
>2>u>�>?R?�?�?   � t   50�0�0%1r1�1�122u2�23�3�34�4�45V5�5�5E6�6�6(7�7(8�8�8%9b9�9�9E:�:�:%;u;�;<U<�<�<F=�=�=5>q>�>�>�>E?�?�?   � x   0e0�01e1�12e2�2�2%3f3�3�3E4�4�45o5�5�56\6�67|78b8h8�8�8�8�8�8�89H9[9u9�9�9�9�9�9�9�9�9:t:�:�:;�>m?}?   � �   �0 1g1�1�1�1�1�12_2�2343�34�4V5�5�5�56;6�7L8t8T9t9�9�9:1:T:�:�:�:;4;d;�;�;M<T<[<b<i<p<w<~<�<�<�<�<�<�<�<�<�<�<�<�<�<�<(=E=y=->�>�?�?�?�?   � D  010G0Y0^0d0j0�0�0�0�0�0�01I1O1j1�1�1�1"2O2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33
33/3B3^3�3J44�4�4�4�4�4�4�45!5(5,5054585<5@5D5�5�5�5�5�566,63686<6@6a6�6�6�6�6�6�6�6�6�6�6*7074787<7�788j8t8�8�8�8919�9�9�9�9�9:�:�:�:�:�:�:];w;�;�;�;P<b<�<�<�<�<�<�<=%=*=>->3><>C>b>�>??&?.?B?M?R?d?n?u?�?�?�?�?�?�?�?�?�?   � d  90>0I0N0l0�0�0.1G1s1y1�1�1�1�1�1�1�1�1�122"262=2W2a2g2s2�2�2�2�2�2�2�2�2�2�2�2�2333<3F3a3�3�3�3�3�3�34�4�4�4�4�4>5Q5W5c5i5x5~5�5�5�5�5�5�5�5�5�5�5�5�5�5�5666!6&6+61656;6@6F6N6Z6p6{6�6�6�6�6�6�6�6�6�6�6�67?7H7T7�7�7�7�7�7�7�7848:8l8�8�899=9V9�9�9�9+:1:S:q:�:�:�:�:�:>;I;Q;c;n;=-=5=;=@=H=�=�=�=�=�=�=>>D>�>�>�>�> ??$?)?�?�?�?�?�?�?�? � \   	000-060B0K0R0\0b0h0�011 1&1�12_2C3K3d3~3�3�344)41494E4i4q4l5t5�5�588�8�8%>�>     |0�0�0�01
11-13191?1E1K1R1Y1`1g1n1u1|1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�122!2)242J2X2{23"333G3[3�3�3�3�3�3�3�30454]44�4�4�4�45*5�7�7�7�7�7�7�7�78&8,858H8l8�89/959<9I9P9V9^9d9p9u9�;�;�;�;�;�;<<<+<><I<O<U<Z<c<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<==&=7===N=�=    �   I1U1�1�1�1-2 444.4I4j4}4�4�4�455{5�5�5�5666(6M6V6_6l6�6�6�6�6�6�6�6�6�6�677L7P7T7X7\7`7d7h7l7p7t7x7|7�7�7T8�8�8�8)9�98:�:k;l<|<�<�<�<�<�<=�=!>1>=>O>_>k>h?�?�?�?�?   D   80`0e7�8�89�9�9�9:a;|;�;q<{<�<�<�<�=�=�=�=�=�=v?{?�?�?�?�? 0 �   .0e0p0z00�0�0�0�0�011c1h1o1t1{1�1�1�1�1�2�2�2�2�2�2�2�2�2	33P3}3B4h4�4�4<5�5�5�56H6�6778�8�8�8�8�8�8979?9I9b9l99�9�9: :�:�:�:W;v;�;�;
<<7<?<G<^<w<�<�<�<�<�<�<�<= =.=�=�=�=�=�=L>>�>"?(?y??�?�?�? @ L    00S0�0�0�13"3+4�4�445L5�5�5�5P898:^:}:<�=�=�=�=�=�=�=�=.>;>n?�? P �   @0
1?1X1_1g1l1p1t1�1�1�1�1�1�1�1�1�1 22N2T2X2\2`2�2�2�2�2�2�2 3!3K3}3�3�3�3�3�3�3�3�3�3�3�3�3�3�5�7�7�8�8�8�8�8�8�8�8�8�8929C9J9Y9^9k9y9�9::~;�;�;�=R?m?�?�?�?   ` p   01x1�1�1M284K4]4�4�4�4�4 5�5r8�8�8�8�8�8�8�899|9�9�9�9�9�9�9�9�9�:	;�;�;�;�;�;�;�;/<_<�<�=�=F>?�?   p �   	00�0�0�01171U1�1�1z2�2�3�3�4�4�4(6�6�7�7�7�78�8�8�8k9�9�9::,:=:H:V:d:k:z:�:�:�:�:�:�:�:;G;Q;Z;};�;�;�;=!=�>�?�? � T   �0p1	22�2�2�2g3~3455�5�6K7Q7�7�7	8�8�8�8{9K<b<w?{??�?�?�?�?�?�?�?�?�?�? � $   �0�0�0�061[1;�>?'?D?n?�?�? � �   �0�0(181S1s1�1�12*2�2�2�2�2�2�2�2�233'323G3N3T3j3�3&4�4�4�4�455"505�5"6-6P6�6�6P9V9[9a9k9z9:~:�:�:	;;r;�;�;�;�;*<Y<�=�=�=�=�=>>+>   �   $1014181<1@1L1P1�1�1�1�1�1�1�1�1�1 22222222 2$2,2024282<2@2D2H2L2�3�3�3�3�3�3�344 4$4(4,4044484<4P4T4X4\4`4d4h4l4p4t4x4|4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4�4 55555555 5$5(5,5054585<5@5D5H5L5P5T5X5\5`5d587<7@7D7H7�7�7�7�7�7�7�7�7 888880949   � �   �5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7,7074787<7@7D7H7L7P7T7 � P  �3�3�3�3�3�3�3�34440444D4H4L4P4X4p4�4�4�4�4�4�4�4�4�4�4�4�4�4�45$5(5<5@5P5T5X5\5d5|5�5�5�5�5�5�5�5�5�5�5666 6$6,6D6T6X6h6l6|6�6�6�6�6�6�6�6�6�6�6�6�6�67$7(787<7@7D7L7d7t7x7�7�7�7�7�7�7�7�7�7�78888$8<8L8P8`8d8h8p8�8�8�8�8�8�8�8�8�8�8�8 99T9X9x9�9�9�9�9:8:D:\:`:�:�:�:�:�:�: ;; ;@;`;�;�;�;�;�;�; < <@<`<�<�<�<�<�<= � �   00 080X0x0�0�0�0�0�0�0�01014181<1@1D1`1x1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1�1242X2t2x2|2�2�2�2�2�2�2�2�2�2�2�2�2�2�2 33333 3 44444444 4$444<4D4L4T4\4d4l4t4|4�4�4�4�4�4�4�4�4�4�4�4�4�488888"8&8*8.82868:8>8B8F8J8N8R8V8Z8^8b8f8j8n8r8v8z8~8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�899
99x9�9�9�9�9�9�9�9�9�9�9 ::0>(?,?L?T?\?d?l?t?|?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   �   0000$0,0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0�0 11111111 1$1(1,101@1H1L1P1T1X1\1`1d1h1l1x1�1�1�4�4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              